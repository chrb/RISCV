-- Copyright (C) 1991-2013 Altera Corporation
-- Your use of Altera Corporation's design tools, logic functions 
-- and other software and tools, and its AMPP partner logic 
-- functions, and any output files from any of the foregoing 
-- (including device programming or simulation files), and any 
-- associated documentation or information are expressly subject 
-- to the terms and conditions of the Altera Program License 
-- Subscription Agreement, Altera MegaCore Function License 
-- Agreement, or other applicable license agreement, including, 
-- without limitation, that your use is for the sole purpose of 
-- programming logic devices manufactured by Altera and sold by 
-- Altera or its authorized distributors.  Please refer to the 
-- applicable agreement for further details.

-- PROGRAM		"Quartus II 32-bit"
-- VERSION		"Version 13.0.1 Build 232 06/12/2013 Service Pack 1 SJ Full Version"
-- CREATED		"Fri Feb  5 11:04:18 2016"

LIBRARY ieee;
USE ieee.std_logic_1164.all; 

LIBRARY work;

ENTITY RISCV_SDRAM IS 
	PORT
	(
		CLOCK_50 :  IN  STD_LOGIC;
		m_waitrequest :  IN  STD_LOGIC;
		m_readdatavalid :  IN  STD_LOGIC;
		KEY :  IN  STD_LOGIC_VECTOR(1 TO 1);
		m_readdata :  IN  STD_LOGIC_VECTOR(31 DOWNTO 0);
		m_write :  OUT  STD_LOGIC;
		m_read :  OUT  STD_LOGIC;
		HEX0 :  OUT  STD_LOGIC_VECTOR(6 DOWNTO 0);
		HEX1 :  OUT  STD_LOGIC_VECTOR(6 DOWNTO 0);
		HEX2 :  OUT  STD_LOGIC_VECTOR(6 DOWNTO 0);
		HEX3 :  OUT  STD_LOGIC_VECTOR(6 DOWNTO 0);
		m_address :  OUT  STD_LOGIC_VECTOR(20 DOWNTO 0);
		m_byteenable :  OUT  STD_LOGIC_VECTOR(3 DOWNTO 0);
		m_writedata :  OUT  STD_LOGIC_VECTOR(31 DOWNTO 0)
	);
END RISCV_SDRAM;

ARCHITECTURE bdf_type OF RISCV_SDRAM IS 

COMPONENT sevenseg
	PORT(Set : IN STD_LOGIC;
		 Clk : IN STD_LOGIC;
		 nRst : IN STD_LOGIC;
		 V : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
		 Hex0 : OUT STD_LOGIC_VECTOR(6 DOWNTO 0);
		 Hex1 : OUT STD_LOGIC_VECTOR(6 DOWNTO 0);
		 Hex2 : OUT STD_LOGIC_VECTOR(6 DOWNTO 0);
		 Hex3 : OUT STD_LOGIC_VECTOR(6 DOWNTO 0)
	);
END COMPONENT;

COMPONENT instrmem
	PORT(clock : IN STD_LOGIC;
		 address : IN STD_LOGIC_VECTOR(9 DOWNTO 0);
		 q : OUT STD_LOGIC_VECTOR(31 DOWNTO 0)
	);
END COMPONENT;

COMPONENT fetchstage
	PORT(StallI : IN STD_LOGIC;
		 Clk : IN STD_LOGIC;
		 nRst : IN STD_LOGIC;
		 PCI : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
		 StallO : OUT STD_LOGIC;
		 PCO : OUT STD_LOGIC_VECTOR(31 DOWNTO 0)
	);
END COMPONENT;

COMPONENT fetch
	PORT(StallI : IN STD_LOGIC;
		 Jump : IN STD_LOGIC;
		 InterlockI : IN STD_LOGIC;
		 JumpTarget : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
		 PCOld : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
		 ImemAddr : OUT STD_LOGIC_VECTOR(9 DOWNTO 0);
		 PCNext : OUT STD_LOGIC_VECTOR(31 DOWNTO 0)
	);
END COMPONENT;

COMPONENT sdraminterface
	PORT(logic_write : IN STD_LOGIC;
		 logic_read : IN STD_LOGIC;
		 logic_StallI : IN STD_LOGIC;
		 m_readdatavalid : IN STD_LOGIC;
		 m_waitrequest : IN STD_LOGIC;
		 Clk : IN STD_LOGIC;
		 nRst : IN STD_LOGIC;
		 logic_address : IN STD_LOGIC_VECTOR(9 DOWNTO 0);
		 logic_byteenable : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
		 logic_writedata : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
		 m_readdata : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
		 logic_StallO : OUT STD_LOGIC;
		 m_write : OUT STD_LOGIC;
		 m_read : OUT STD_LOGIC;
		 logic_readdata : OUT STD_LOGIC_VECTOR(31 DOWNTO 0);
		 m_address : OUT STD_LOGIC_VECTOR(20 DOWNTO 0);
		 m_byteenable : OUT STD_LOGIC_VECTOR(3 DOWNTO 0);
		 m_writedata : OUT STD_LOGIC_VECTOR(31 DOWNTO 0)
	);
END COMPONENT;

COMPONENT memmux
	PORT(S : IN STD_LOGIC;
		 A : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
		 B : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
		 FunctI : IN STD_LOGIC_VECTOR(2 DOWNTO 0);
		 MemAddrLowI : IN STD_LOGIC_VECTOR(1 DOWNTO 0);
		 O : OUT STD_LOGIC_VECTOR(31 DOWNTO 0)
	);
END COMPONENT;

COMPONENT decode
	PORT(ClearI : IN STD_LOGIC;
		 InterlockI : IN STD_LOGIC;
		 StallI : IN STD_LOGIC;
		 Insn : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
		 PCNextI : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
		 SelSrc2 : OUT STD_LOGIC;
		 Aux : OUT STD_LOGIC;
		 Jump : OUT STD_LOGIC;
		 JumpRel : OUT STD_LOGIC;
		 MemAccess : OUT STD_LOGIC;
		 MemWrEn : OUT STD_LOGIC;
		 MemRdEn : OUT STD_LOGIC;
		 DestWrEn : OUT STD_LOGIC;
		 SetSevenSegO : OUT STD_LOGIC;
		 InterlockO : OUT STD_LOGIC;
		 StallO : OUT STD_LOGIC;
		 DestRegNo : OUT STD_LOGIC_VECTOR(4 DOWNTO 0);
		 Funct : OUT STD_LOGIC_VECTOR(2 DOWNTO 0);
		 Imm : OUT STD_LOGIC_VECTOR(31 DOWNTO 0);
		 JumpTarget : OUT STD_LOGIC_VECTOR(31 DOWNTO 0);
		 PCNextO : OUT STD_LOGIC_VECTOR(31 DOWNTO 0);
		 SrcRegNo1 : OUT STD_LOGIC_VECTOR(4 DOWNTO 0);
		 SrcRegNo2 : OUT STD_LOGIC_VECTOR(4 DOWNTO 0)
	);
END COMPONENT;

COMPONENT alu
	PORT(Aux : IN STD_LOGIC;
		 JumpI : IN STD_LOGIC;
		 JumpRel : IN STD_LOGIC;
		 MemAccessI : IN STD_LOGIC;
		 MemWrEnI : IN STD_LOGIC;
		 MemRdEnI : IN STD_LOGIC;
		 DestWrEnI : IN STD_LOGIC;
		 ClearI : IN STD_LOGIC;
		 A : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
		 B : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
		 DestRegNoI : IN STD_LOGIC_VECTOR(4 DOWNTO 0);
		 FunctI : IN STD_LOGIC_VECTOR(2 DOWNTO 0);
		 JumpTargetI : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
		 MemWrDataI : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
		 PCNextI : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
		 DestWrEnO : OUT STD_LOGIC;
		 MemAccessO : OUT STD_LOGIC;
		 MemWrEnO : OUT STD_LOGIC;
		 MemRdEnO : OUT STD_LOGIC;
		 JumpO : OUT STD_LOGIC;
		 DestRegNoO : OUT STD_LOGIC_VECTOR(4 DOWNTO 0);
		 FunctO : OUT STD_LOGIC_VECTOR(2 DOWNTO 0);
		 JumpTargetO : OUT STD_LOGIC_VECTOR(31 DOWNTO 0);
		 MemAddr : OUT STD_LOGIC_VECTOR(9 DOWNTO 0);
		 MemAddrLow : OUT STD_LOGIC_VECTOR(1 DOWNTO 0);
		 MemByteEna : OUT STD_LOGIC_VECTOR(3 DOWNTO 0);
		 MemWrDataO : OUT STD_LOGIC_VECTOR(31 DOWNTO 0);
		 X : OUT STD_LOGIC_VECTOR(31 DOWNTO 0)
	);
END COMPONENT;

COMPONENT memstage
	PORT(DestWrEnI : IN STD_LOGIC;
		 MemAccessI : IN STD_LOGIC;
		 Clk : IN STD_LOGIC;
		 nRst : IN STD_LOGIC;
		 DestRegNoI : IN STD_LOGIC_VECTOR(4 DOWNTO 0);
		 DestWrDataI : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
		 FunctI : IN STD_LOGIC_VECTOR(2 DOWNTO 0);
		 MemAddrLowI : IN STD_LOGIC_VECTOR(1 DOWNTO 0);
		 DestWrEnO : OUT STD_LOGIC;
		 MemAccessO : OUT STD_LOGIC;
		 DestRegNoO : OUT STD_LOGIC_VECTOR(4 DOWNTO 0);
		 DestWrDataO : OUT STD_LOGIC_VECTOR(31 DOWNTO 0);
		 FunctO : OUT STD_LOGIC_VECTOR(2 DOWNTO 0);
		 MemAddrLowO : OUT STD_LOGIC_VECTOR(1 DOWNTO 0)
	);
END COMPONENT;

COMPONENT forward
	PORT(ExDestWrEn : IN STD_LOGIC;
		 MemDestWrEn : IN STD_LOGIC;
		 ExDestData : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
		 ExDestRegNo : IN STD_LOGIC_VECTOR(4 DOWNTO 0);
		 MemDestData : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
		 MemDestRegNo : IN STD_LOGIC_VECTOR(4 DOWNTO 0);
		 SrcData1 : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
		 SrcData2 : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
		 SrcRegNo1 : IN STD_LOGIC_VECTOR(4 DOWNTO 0);
		 SrcRegNo2 : IN STD_LOGIC_VECTOR(4 DOWNTO 0);
		 FwdData1 : OUT STD_LOGIC_VECTOR(31 DOWNTO 0);
		 FwdData2 : OUT STD_LOGIC_VECTOR(31 DOWNTO 0)
	);
END COMPONENT;

COMPONENT decodestage
	PORT(ClearI : IN STD_LOGIC;
		 InterlockI : IN STD_LOGIC;
		 StallI : IN STD_LOGIC;
		 Clk : IN STD_LOGIC;
		 nRst : IN STD_LOGIC;
		 InsnI : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
		 PCNextI : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
		 ClearO : OUT STD_LOGIC;
		 InterlockO : OUT STD_LOGIC;
		 StallO : OUT STD_LOGIC;
		 InsnO : OUT STD_LOGIC_VECTOR(31 DOWNTO 0);
		 PCNextO : OUT STD_LOGIC_VECTOR(31 DOWNTO 0)
	);
END COMPONENT;

COMPONENT executestage
	PORT(SelSrc2I : IN STD_LOGIC;
		 AuxI : IN STD_LOGIC;
		 JumpI : IN STD_LOGIC;
		 JumpRelI : IN STD_LOGIC;
		 MemAccessI : IN STD_LOGIC;
		 MemWrEnI : IN STD_LOGIC;
		 MemRdEnI : IN STD_LOGIC;
		 DestWrEnI : IN STD_LOGIC;
		 SetSevenSegI : IN STD_LOGIC;
		 ClearI : IN STD_LOGIC;
		 Clk : IN STD_LOGIC;
		 nRst : IN STD_LOGIC;
		 DestRegNoI : IN STD_LOGIC_VECTOR(4 DOWNTO 0);
		 FunctI : IN STD_LOGIC_VECTOR(2 DOWNTO 0);
		 ImmI : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
		 JumpTargetI : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
		 PCNextI : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
		 SrcData1I : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
		 SrcData2I : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
		 SelSrc2O : OUT STD_LOGIC;
		 AuxO : OUT STD_LOGIC;
		 JumpO : OUT STD_LOGIC;
		 JumpRelO : OUT STD_LOGIC;
		 MemAccessO : OUT STD_LOGIC;
		 MemWrEnO : OUT STD_LOGIC;
		 MemRdEnO : OUT STD_LOGIC;
		 DestWrEnO : OUT STD_LOGIC;
		 ClearO : OUT STD_LOGIC;
		 SetSevenSegO : OUT STD_LOGIC;
		 DestRegNoO : OUT STD_LOGIC_VECTOR(4 DOWNTO 0);
		 FunctO : OUT STD_LOGIC_VECTOR(2 DOWNTO 0);
		 ImmO : OUT STD_LOGIC_VECTOR(31 DOWNTO 0);
		 JumpTargetO : OUT STD_LOGIC_VECTOR(31 DOWNTO 0);
		 PCNextO : OUT STD_LOGIC_VECTOR(31 DOWNTO 0);
		 SrcData1O : OUT STD_LOGIC_VECTOR(31 DOWNTO 0);
		 SrcData2O : OUT STD_LOGIC_VECTOR(31 DOWNTO 0)
	);
END COMPONENT;

COMPONENT regset
	PORT(WrEn : IN STD_LOGIC;
		 Clk : IN STD_LOGIC;
		 nRst : IN STD_LOGIC;
		 RdRegNo1 : IN STD_LOGIC_VECTOR(4 DOWNTO 0);
		 RdRegNo2 : IN STD_LOGIC_VECTOR(4 DOWNTO 0);
		 WrData : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
		 WrRegNo : IN STD_LOGIC_VECTOR(4 DOWNTO 0);
		 RdData1 : OUT STD_LOGIC_VECTOR(31 DOWNTO 0);
		 RdData2 : OUT STD_LOGIC_VECTOR(31 DOWNTO 0)
	);
END COMPONENT;

COMPONENT mux32bit
	PORT(S : IN STD_LOGIC;
		 A : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
		 B : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
		 O : OUT STD_LOGIC_VECTOR(31 DOWNTO 0)
	);
END COMPONENT;

SIGNAL	SYNTHESIZED_WIRE_0 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_87 :  STD_LOGIC_VECTOR(31 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_2 :  STD_LOGIC_VECTOR(9 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_88 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_89 :  STD_LOGIC_VECTOR(31 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_5 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_90 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_91 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_8 :  STD_LOGIC_VECTOR(31 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_9 :  STD_LOGIC_VECTOR(31 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_10 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_11 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_12 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_13 :  STD_LOGIC_VECTOR(9 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_14 :  STD_LOGIC_VECTOR(3 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_15 :  STD_LOGIC_VECTOR(31 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_16 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_17 :  STD_LOGIC_VECTOR(31 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_18 :  STD_LOGIC_VECTOR(31 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_19 :  STD_LOGIC_VECTOR(2 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_20 :  STD_LOGIC_VECTOR(1 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_21 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_22 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_23 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_24 :  STD_LOGIC_VECTOR(31 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_25 :  STD_LOGIC_VECTOR(31 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_26 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_27 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_28 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_29 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_30 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_31 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_92 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_33 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_35 :  STD_LOGIC_VECTOR(31 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_93 :  STD_LOGIC_VECTOR(4 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_37 :  STD_LOGIC_VECTOR(2 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_38 :  STD_LOGIC_VECTOR(31 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_94 :  STD_LOGIC_VECTOR(31 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_40 :  STD_LOGIC_VECTOR(31 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_41 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_42 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_43 :  STD_LOGIC_VECTOR(4 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_95 :  STD_LOGIC_VECTOR(31 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_45 :  STD_LOGIC_VECTOR(2 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_46 :  STD_LOGIC_VECTOR(1 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_96 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_97 :  STD_LOGIC_VECTOR(31 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_98 :  STD_LOGIC_VECTOR(4 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_53 :  STD_LOGIC_VECTOR(31 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_54 :  STD_LOGIC_VECTOR(31 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_99 :  STD_LOGIC_VECTOR(4 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_100 :  STD_LOGIC_VECTOR(4 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_60 :  STD_LOGIC_VECTOR(31 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_62 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_63 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_64 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_65 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_66 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_67 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_68 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_69 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_70 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_72 :  STD_LOGIC_VECTOR(4 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_73 :  STD_LOGIC_VECTOR(2 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_74 :  STD_LOGIC_VECTOR(31 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_75 :  STD_LOGIC_VECTOR(31 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_76 :  STD_LOGIC_VECTOR(31 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_77 :  STD_LOGIC_VECTOR(31 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_78 :  STD_LOGIC_VECTOR(31 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_84 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_86 :  STD_LOGIC_VECTOR(31 DOWNTO 0);


BEGIN 



b2v_inst : sevenseg
PORT MAP(Set => SYNTHESIZED_WIRE_0,
		 Clk => CLOCK_50,
		 nRst => KEY(1),
		 V => SYNTHESIZED_WIRE_87,
		 Hex0 => HEX0,
		 Hex1 => HEX1,
		 Hex2 => HEX2,
		 Hex3 => HEX3);


b2v_inst1 : instrmem
PORT MAP(clock => CLOCK_50,
		 address => SYNTHESIZED_WIRE_2,
		 q => SYNTHESIZED_WIRE_60);


b2v_inst10 : fetchstage
PORT MAP(StallI => SYNTHESIZED_WIRE_88,
		 Clk => CLOCK_50,
		 nRst => KEY(1),
		 PCI => SYNTHESIZED_WIRE_89,
		 StallO => SYNTHESIZED_WIRE_5,
		 PCO => SYNTHESIZED_WIRE_9);


b2v_inst11 : fetch
PORT MAP(StallI => SYNTHESIZED_WIRE_5,
		 Jump => SYNTHESIZED_WIRE_90,
		 InterlockI => SYNTHESIZED_WIRE_91,
		 JumpTarget => SYNTHESIZED_WIRE_8,
		 PCOld => SYNTHESIZED_WIRE_9,
		 ImemAddr => SYNTHESIZED_WIRE_2,
		 PCNext => SYNTHESIZED_WIRE_89);


b2v_inst12 : sdraminterface
PORT MAP(logic_write => SYNTHESIZED_WIRE_10,
		 logic_read => SYNTHESIZED_WIRE_11,
		 logic_StallI => SYNTHESIZED_WIRE_12,
		 m_readdatavalid => m_readdatavalid,
		 m_waitrequest => m_waitrequest,
		 Clk => CLOCK_50,
		 nRst => KEY(1),
		 logic_address => SYNTHESIZED_WIRE_13,
		 logic_byteenable => SYNTHESIZED_WIRE_14,
		 logic_writedata => SYNTHESIZED_WIRE_15,
		 m_readdata => m_readdata,
		 logic_StallO => SYNTHESIZED_WIRE_88,
		 m_write => m_write,
		 m_read => m_read,
		 logic_readdata => SYNTHESIZED_WIRE_18,
		 m_address => m_address,
		 m_byteenable => m_byteenable,
		 m_writedata => m_writedata);


b2v_inst17 : memmux
PORT MAP(S => SYNTHESIZED_WIRE_16,
		 A => SYNTHESIZED_WIRE_17,
		 B => SYNTHESIZED_WIRE_18,
		 FunctI => SYNTHESIZED_WIRE_19,
		 MemAddrLowI => SYNTHESIZED_WIRE_20,
		 O => SYNTHESIZED_WIRE_97);


b2v_inst2 : decode
PORT MAP(ClearI => SYNTHESIZED_WIRE_21,
		 InterlockI => SYNTHESIZED_WIRE_22,
		 StallI => SYNTHESIZED_WIRE_23,
		 Insn => SYNTHESIZED_WIRE_24,
		 PCNextI => SYNTHESIZED_WIRE_25,
		 SelSrc2 => SYNTHESIZED_WIRE_62,
		 Aux => SYNTHESIZED_WIRE_63,
		 Jump => SYNTHESIZED_WIRE_64,
		 JumpRel => SYNTHESIZED_WIRE_65,
		 MemAccess => SYNTHESIZED_WIRE_66,
		 MemWrEn => SYNTHESIZED_WIRE_67,
		 MemRdEn => SYNTHESIZED_WIRE_68,
		 DestWrEn => SYNTHESIZED_WIRE_69,
		 SetSevenSegO => SYNTHESIZED_WIRE_70,
		 InterlockO => SYNTHESIZED_WIRE_91,
		 StallO => SYNTHESIZED_WIRE_12,
		 DestRegNo => SYNTHESIZED_WIRE_72,
		 Funct => SYNTHESIZED_WIRE_73,
		 Imm => SYNTHESIZED_WIRE_74,
		 JumpTarget => SYNTHESIZED_WIRE_75,
		 PCNextO => SYNTHESIZED_WIRE_76,
		 SrcRegNo1 => SYNTHESIZED_WIRE_99,
		 SrcRegNo2 => SYNTHESIZED_WIRE_100);


b2v_inst3 : alu
PORT MAP(Aux => SYNTHESIZED_WIRE_26,
		 JumpI => SYNTHESIZED_WIRE_27,
		 JumpRel => SYNTHESIZED_WIRE_28,
		 MemAccessI => SYNTHESIZED_WIRE_29,
		 MemWrEnI => SYNTHESIZED_WIRE_30,
		 MemRdEnI => SYNTHESIZED_WIRE_31,
		 DestWrEnI => SYNTHESIZED_WIRE_92,
		 ClearI => SYNTHESIZED_WIRE_33,
		 A => SYNTHESIZED_WIRE_87,
		 B => SYNTHESIZED_WIRE_35,
		 DestRegNoI => SYNTHESIZED_WIRE_93,
		 FunctI => SYNTHESIZED_WIRE_37,
		 JumpTargetI => SYNTHESIZED_WIRE_38,
		 MemWrDataI => SYNTHESIZED_WIRE_94,
		 PCNextI => SYNTHESIZED_WIRE_40,
		 DestWrEnO => SYNTHESIZED_WIRE_41,
		 MemAccessO => SYNTHESIZED_WIRE_42,
		 MemWrEnO => SYNTHESIZED_WIRE_10,
		 MemRdEnO => SYNTHESIZED_WIRE_11,
		 JumpO => SYNTHESIZED_WIRE_90,
		 DestRegNoO => SYNTHESIZED_WIRE_43,
		 FunctO => SYNTHESIZED_WIRE_45,
		 JumpTargetO => SYNTHESIZED_WIRE_8,
		 MemAddr => SYNTHESIZED_WIRE_13,
		 MemAddrLow => SYNTHESIZED_WIRE_46,
		 MemByteEna => SYNTHESIZED_WIRE_14,
		 MemWrDataO => SYNTHESIZED_WIRE_15,
		 X => SYNTHESIZED_WIRE_95);


b2v_inst4 : memstage
PORT MAP(DestWrEnI => SYNTHESIZED_WIRE_41,
		 MemAccessI => SYNTHESIZED_WIRE_42,
		 Clk => CLOCK_50,
		 nRst => KEY(1),
		 DestRegNoI => SYNTHESIZED_WIRE_43,
		 DestWrDataI => SYNTHESIZED_WIRE_95,
		 FunctI => SYNTHESIZED_WIRE_45,
		 MemAddrLowI => SYNTHESIZED_WIRE_46,
		 DestWrEnO => SYNTHESIZED_WIRE_96,
		 MemAccessO => SYNTHESIZED_WIRE_16,
		 DestRegNoO => SYNTHESIZED_WIRE_98,
		 DestWrDataO => SYNTHESIZED_WIRE_17,
		 FunctO => SYNTHESIZED_WIRE_19,
		 MemAddrLowO => SYNTHESIZED_WIRE_20);


b2v_inst5 : forward
PORT MAP(ExDestWrEn => SYNTHESIZED_WIRE_92,
		 MemDestWrEn => SYNTHESIZED_WIRE_96,
		 ExDestData => SYNTHESIZED_WIRE_95,
		 ExDestRegNo => SYNTHESIZED_WIRE_93,
		 MemDestData => SYNTHESIZED_WIRE_97,
		 MemDestRegNo => SYNTHESIZED_WIRE_98,
		 SrcData1 => SYNTHESIZED_WIRE_53,
		 SrcData2 => SYNTHESIZED_WIRE_54,
		 SrcRegNo1 => SYNTHESIZED_WIRE_99,
		 SrcRegNo2 => SYNTHESIZED_WIRE_100,
		 FwdData1 => SYNTHESIZED_WIRE_77,
		 FwdData2 => SYNTHESIZED_WIRE_78);


b2v_inst6 : decodestage
PORT MAP(ClearI => SYNTHESIZED_WIRE_90,
		 InterlockI => SYNTHESIZED_WIRE_91,
		 StallI => SYNTHESIZED_WIRE_88,
		 Clk => CLOCK_50,
		 nRst => KEY(1),
		 InsnI => SYNTHESIZED_WIRE_60,
		 PCNextI => SYNTHESIZED_WIRE_89,
		 ClearO => SYNTHESIZED_WIRE_21,
		 InterlockO => SYNTHESIZED_WIRE_22,
		 StallO => SYNTHESIZED_WIRE_23,
		 InsnO => SYNTHESIZED_WIRE_24,
		 PCNextO => SYNTHESIZED_WIRE_25);


b2v_inst7 : executestage
PORT MAP(SelSrc2I => SYNTHESIZED_WIRE_62,
		 AuxI => SYNTHESIZED_WIRE_63,
		 JumpI => SYNTHESIZED_WIRE_64,
		 JumpRelI => SYNTHESIZED_WIRE_65,
		 MemAccessI => SYNTHESIZED_WIRE_66,
		 MemWrEnI => SYNTHESIZED_WIRE_67,
		 MemRdEnI => SYNTHESIZED_WIRE_68,
		 DestWrEnI => SYNTHESIZED_WIRE_69,
		 SetSevenSegI => SYNTHESIZED_WIRE_70,
		 ClearI => SYNTHESIZED_WIRE_90,
		 Clk => CLOCK_50,
		 nRst => KEY(1),
		 DestRegNoI => SYNTHESIZED_WIRE_72,
		 FunctI => SYNTHESIZED_WIRE_73,
		 ImmI => SYNTHESIZED_WIRE_74,
		 JumpTargetI => SYNTHESIZED_WIRE_75,
		 PCNextI => SYNTHESIZED_WIRE_76,
		 SrcData1I => SYNTHESIZED_WIRE_77,
		 SrcData2I => SYNTHESIZED_WIRE_78,
		 SelSrc2O => SYNTHESIZED_WIRE_84,
		 AuxO => SYNTHESIZED_WIRE_26,
		 JumpO => SYNTHESIZED_WIRE_27,
		 JumpRelO => SYNTHESIZED_WIRE_28,
		 MemAccessO => SYNTHESIZED_WIRE_29,
		 MemWrEnO => SYNTHESIZED_WIRE_30,
		 MemRdEnO => SYNTHESIZED_WIRE_31,
		 DestWrEnO => SYNTHESIZED_WIRE_92,
		 ClearO => SYNTHESIZED_WIRE_33,
		 SetSevenSegO => SYNTHESIZED_WIRE_0,
		 DestRegNoO => SYNTHESIZED_WIRE_93,
		 FunctO => SYNTHESIZED_WIRE_37,
		 ImmO => SYNTHESIZED_WIRE_86,
		 JumpTargetO => SYNTHESIZED_WIRE_38,
		 PCNextO => SYNTHESIZED_WIRE_40,
		 SrcData1O => SYNTHESIZED_WIRE_87,
		 SrcData2O => SYNTHESIZED_WIRE_94);


b2v_inst8 : regset
PORT MAP(WrEn => SYNTHESIZED_WIRE_96,
		 Clk => CLOCK_50,
		 nRst => KEY(1),
		 RdRegNo1 => SYNTHESIZED_WIRE_99,
		 RdRegNo2 => SYNTHESIZED_WIRE_100,
		 WrData => SYNTHESIZED_WIRE_97,
		 WrRegNo => SYNTHESIZED_WIRE_98,
		 RdData1 => SYNTHESIZED_WIRE_53,
		 RdData2 => SYNTHESIZED_WIRE_54);


b2v_inst9 : mux32bit
PORT MAP(S => SYNTHESIZED_WIRE_84,
		 A => SYNTHESIZED_WIRE_94,
		 B => SYNTHESIZED_WIRE_86,
		 O => SYNTHESIZED_WIRE_35);


END bdf_type;