-- SDRAM.vhd

-- Generated using ACDS version 13.0sp1 232 at 2016.02.05.11:39:02

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity SDRAM is
	port (
		clk_clk       : in std_logic := '0'; --   clk.clk
		reset_reset_n : in std_logic := '0'  -- reset.reset_n
	);
end entity SDRAM;

architecture rtl of SDRAM is
	component SDRAM_sdram_controller is
		port (
			clk            : in    std_logic                     := 'X';             -- clk
			reset_n        : in    std_logic                     := 'X';             -- reset_n
			az_addr        : in    std_logic_vector(20 downto 0) := (others => 'X'); -- address
			az_be_n        : in    std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable_n
			az_cs          : in    std_logic                     := 'X';             -- chipselect
			az_data        : in    std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			az_rd_n        : in    std_logic                     := 'X';             -- read_n
			az_wr_n        : in    std_logic                     := 'X';             -- write_n
			za_data        : out   std_logic_vector(31 downto 0);                    -- readdata
			za_valid       : out   std_logic;                                        -- readdatavalid
			za_waitrequest : out   std_logic;                                        -- waitrequest
			zs_addr        : out   std_logic_vector(10 downto 0);                    -- export
			zs_ba          : out   std_logic_vector(1 downto 0);                     -- export
			zs_cas_n       : out   std_logic;                                        -- export
			zs_cke         : out   std_logic;                                        -- export
			zs_cs_n        : out   std_logic;                                        -- export
			zs_dq          : inout std_logic_vector(31 downto 0) := (others => 'X'); -- export
			zs_dqm         : out   std_logic_vector(3 downto 0);                     -- export
			zs_ras_n       : out   std_logic;                                        -- export
			zs_we_n        : out   std_logic                                         -- export
		);
	end component SDRAM_sdram_controller;

	component SDRAM_SDRAM_Master is
		port (
			CLOCK_50        : in  std_logic                     := 'X';             -- clk
			KEY             : in  std_logic                     := 'X';             -- reset
			HEX0            : out std_logic_vector(6 downto 0);                     -- export
			HEX1            : out std_logic_vector(6 downto 0);                     -- export
			HEX3            : out std_logic_vector(6 downto 0);                     -- export
			HEX2            : out std_logic_vector(6 downto 0);                     -- export
			m_waitrequest   : in  std_logic                     := 'X';             -- waitrequest
			m_readdatavalid : in  std_logic                     := 'X';             -- readdatavalid
			m_readdata      : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			m_write         : out std_logic;                                        -- write
			m_read          : out std_logic;                                        -- read
			m_address       : out std_logic_vector(20 downto 0);                    -- address
			m_byteenable    : out std_logic_vector(3 downto 0);                     -- byteenable
			m_writedata     : out std_logic_vector(31 downto 0)                     -- writedata
		);
	end component SDRAM_SDRAM_Master;

	component altera_merlin_master_translator is
		generic (
			AV_ADDRESS_W                : integer := 32;
			AV_DATA_W                   : integer := 32;
			AV_BURSTCOUNT_W             : integer := 4;
			AV_BYTEENABLE_W             : integer := 4;
			UAV_ADDRESS_W               : integer := 38;
			UAV_BURSTCOUNT_W            : integer := 10;
			USE_READ                    : integer := 1;
			USE_WRITE                   : integer := 1;
			USE_BEGINBURSTTRANSFER      : integer := 0;
			USE_BEGINTRANSFER           : integer := 0;
			USE_CHIPSELECT              : integer := 0;
			USE_BURSTCOUNT              : integer := 1;
			USE_READDATAVALID           : integer := 1;
			USE_WAITREQUEST             : integer := 1;
			USE_READRESPONSE            : integer := 0;
			USE_WRITERESPONSE           : integer := 0;
			AV_SYMBOLS_PER_WORD         : integer := 4;
			AV_ADDRESS_SYMBOLS          : integer := 0;
			AV_BURSTCOUNT_SYMBOLS       : integer := 0;
			AV_CONSTANT_BURST_BEHAVIOR  : integer := 0;
			UAV_CONSTANT_BURST_BEHAVIOR : integer := 0;
			AV_LINEWRAPBURSTS           : integer := 0;
			AV_REGISTERINCOMINGSIGNALS  : integer := 0
		);
		port (
			clk                      : in  std_logic                     := 'X';             -- clk
			reset                    : in  std_logic                     := 'X';             -- reset
			uav_address              : out std_logic_vector(22 downto 0);                    -- address
			uav_burstcount           : out std_logic_vector(2 downto 0);                     -- burstcount
			uav_read                 : out std_logic;                                        -- read
			uav_write                : out std_logic;                                        -- write
			uav_waitrequest          : in  std_logic                     := 'X';             -- waitrequest
			uav_readdatavalid        : in  std_logic                     := 'X';             -- readdatavalid
			uav_byteenable           : out std_logic_vector(3 downto 0);                     -- byteenable
			uav_readdata             : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			uav_writedata            : out std_logic_vector(31 downto 0);                    -- writedata
			uav_lock                 : out std_logic;                                        -- lock
			uav_debugaccess          : out std_logic;                                        -- debugaccess
			av_address               : in  std_logic_vector(20 downto 0) := (others => 'X'); -- address
			av_waitrequest           : out std_logic;                                        -- waitrequest
			av_byteenable            : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			av_read                  : in  std_logic                     := 'X';             -- read
			av_readdata              : out std_logic_vector(31 downto 0);                    -- readdata
			av_readdatavalid         : out std_logic;                                        -- readdatavalid
			av_write                 : in  std_logic                     := 'X';             -- write
			av_writedata             : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			av_burstcount            : in  std_logic_vector(0 downto 0)  := (others => 'X'); -- burstcount
			av_beginbursttransfer    : in  std_logic                     := 'X';             -- beginbursttransfer
			av_begintransfer         : in  std_logic                     := 'X';             -- begintransfer
			av_chipselect            : in  std_logic                     := 'X';             -- chipselect
			av_lock                  : in  std_logic                     := 'X';             -- lock
			av_debugaccess           : in  std_logic                     := 'X';             -- debugaccess
			uav_clken                : out std_logic;                                        -- clken
			av_clken                 : in  std_logic                     := 'X';             -- clken
			uav_response             : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- response
			av_response              : out std_logic_vector(1 downto 0);                     -- response
			uav_writeresponserequest : out std_logic;                                        -- writeresponserequest
			uav_writeresponsevalid   : in  std_logic                     := 'X';             -- writeresponsevalid
			av_writeresponserequest  : in  std_logic                     := 'X';             -- writeresponserequest
			av_writeresponsevalid    : out std_logic                                         -- writeresponsevalid
		);
	end component altera_merlin_master_translator;

	component altera_merlin_slave_translator is
		generic (
			AV_ADDRESS_W                   : integer := 30;
			AV_DATA_W                      : integer := 32;
			UAV_DATA_W                     : integer := 32;
			AV_BURSTCOUNT_W                : integer := 4;
			AV_BYTEENABLE_W                : integer := 4;
			UAV_BYTEENABLE_W               : integer := 4;
			UAV_ADDRESS_W                  : integer := 32;
			UAV_BURSTCOUNT_W               : integer := 4;
			AV_READLATENCY                 : integer := 0;
			USE_READDATAVALID              : integer := 1;
			USE_WAITREQUEST                : integer := 1;
			USE_UAV_CLKEN                  : integer := 0;
			USE_READRESPONSE               : integer := 0;
			USE_WRITERESPONSE              : integer := 0;
			AV_SYMBOLS_PER_WORD            : integer := 4;
			AV_ADDRESS_SYMBOLS             : integer := 0;
			AV_BURSTCOUNT_SYMBOLS          : integer := 0;
			AV_CONSTANT_BURST_BEHAVIOR     : integer := 0;
			UAV_CONSTANT_BURST_BEHAVIOR    : integer := 0;
			AV_REQUIRE_UNALIGNED_ADDRESSES : integer := 0;
			CHIPSELECT_THROUGH_READLATENCY : integer := 0;
			AV_READ_WAIT_CYCLES            : integer := 0;
			AV_WRITE_WAIT_CYCLES           : integer := 0;
			AV_SETUP_WAIT_CYCLES           : integer := 0;
			AV_DATA_HOLD_CYCLES            : integer := 0
		);
		port (
			clk                      : in  std_logic                     := 'X';             -- clk
			reset                    : in  std_logic                     := 'X';             -- reset
			uav_address              : in  std_logic_vector(22 downto 0) := (others => 'X'); -- address
			uav_burstcount           : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- burstcount
			uav_read                 : in  std_logic                     := 'X';             -- read
			uav_write                : in  std_logic                     := 'X';             -- write
			uav_waitrequest          : out std_logic;                                        -- waitrequest
			uav_readdatavalid        : out std_logic;                                        -- readdatavalid
			uav_byteenable           : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			uav_readdata             : out std_logic_vector(31 downto 0);                    -- readdata
			uav_writedata            : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			uav_lock                 : in  std_logic                     := 'X';             -- lock
			uav_debugaccess          : in  std_logic                     := 'X';             -- debugaccess
			av_address               : out std_logic_vector(20 downto 0);                    -- address
			av_write                 : out std_logic;                                        -- write
			av_read                  : out std_logic;                                        -- read
			av_readdata              : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			av_writedata             : out std_logic_vector(31 downto 0);                    -- writedata
			av_byteenable            : out std_logic_vector(3 downto 0);                     -- byteenable
			av_readdatavalid         : in  std_logic                     := 'X';             -- readdatavalid
			av_waitrequest           : in  std_logic                     := 'X';             -- waitrequest
			av_chipselect            : out std_logic;                                        -- chipselect
			av_begintransfer         : out std_logic;                                        -- begintransfer
			av_beginbursttransfer    : out std_logic;                                        -- beginbursttransfer
			av_burstcount            : out std_logic_vector(0 downto 0);                     -- burstcount
			av_writebyteenable       : out std_logic_vector(3 downto 0);                     -- writebyteenable
			av_lock                  : out std_logic;                                        -- lock
			av_clken                 : out std_logic;                                        -- clken
			uav_clken                : in  std_logic                     := 'X';             -- clken
			av_debugaccess           : out std_logic;                                        -- debugaccess
			av_outputenable          : out std_logic;                                        -- outputenable
			uav_response             : out std_logic_vector(1 downto 0);                     -- response
			av_response              : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- response
			uav_writeresponserequest : in  std_logic                     := 'X';             -- writeresponserequest
			uav_writeresponsevalid   : out std_logic;                                        -- writeresponsevalid
			av_writeresponserequest  : out std_logic;                                        -- writeresponserequest
			av_writeresponsevalid    : in  std_logic                     := 'X'              -- writeresponsevalid
		);
	end component altera_merlin_slave_translator;

	component altera_reset_controller is
		generic (
			NUM_RESET_INPUTS        : integer := 6;
			OUTPUT_RESET_SYNC_EDGES : string  := "deassert";
			SYNC_DEPTH              : integer := 2;
			RESET_REQUEST_PRESENT   : integer := 0
		);
		port (
			reset_in0  : in  std_logic := 'X'; -- reset
			clk        : in  std_logic := 'X'; -- clk
			reset_out  : out std_logic;        -- reset
			reset_req  : out std_logic;        -- reset_req
			reset_in1  : in  std_logic := 'X'; -- reset
			reset_in2  : in  std_logic := 'X'; -- reset
			reset_in3  : in  std_logic := 'X'; -- reset
			reset_in4  : in  std_logic := 'X'; -- reset
			reset_in5  : in  std_logic := 'X'; -- reset
			reset_in6  : in  std_logic := 'X'; -- reset
			reset_in7  : in  std_logic := 'X'; -- reset
			reset_in8  : in  std_logic := 'X'; -- reset
			reset_in9  : in  std_logic := 'X'; -- reset
			reset_in10 : in  std_logic := 'X'; -- reset
			reset_in11 : in  std_logic := 'X'; -- reset
			reset_in12 : in  std_logic := 'X'; -- reset
			reset_in13 : in  std_logic := 'X'; -- reset
			reset_in14 : in  std_logic := 'X'; -- reset
			reset_in15 : in  std_logic := 'X'  -- reset
		);
	end component altera_reset_controller;

	signal sdram_master_avalon_master_waitrequest                                        : std_logic;                     -- SDRAM_Master_avalon_master_translator:av_waitrequest -> SDRAM_Master:m_waitrequest
	signal sdram_master_avalon_master_writedata                                          : std_logic_vector(31 downto 0); -- SDRAM_Master:m_writedata -> SDRAM_Master_avalon_master_translator:av_writedata
	signal sdram_master_avalon_master_address                                            : std_logic_vector(20 downto 0); -- SDRAM_Master:m_address -> SDRAM_Master_avalon_master_translator:av_address
	signal sdram_master_avalon_master_write                                              : std_logic;                     -- SDRAM_Master:m_write -> SDRAM_Master_avalon_master_translator:av_write
	signal sdram_master_avalon_master_read                                               : std_logic;                     -- SDRAM_Master:m_read -> SDRAM_Master_avalon_master_translator:av_read
	signal sdram_master_avalon_master_readdata                                           : std_logic_vector(31 downto 0); -- SDRAM_Master_avalon_master_translator:av_readdata -> SDRAM_Master:m_readdata
	signal sdram_master_avalon_master_byteenable                                         : std_logic_vector(3 downto 0);  -- SDRAM_Master:m_byteenable -> SDRAM_Master_avalon_master_translator:av_byteenable
	signal sdram_master_avalon_master_readdatavalid                                      : std_logic;                     -- SDRAM_Master_avalon_master_translator:av_readdatavalid -> SDRAM_Master:m_readdatavalid
	signal sdram_master_avalon_master_translator_avalon_universal_master_0_waitrequest   : std_logic;                     -- sdram_controller_s1_translator:uav_waitrequest -> SDRAM_Master_avalon_master_translator:uav_waitrequest
	signal sdram_master_avalon_master_translator_avalon_universal_master_0_burstcount    : std_logic_vector(2 downto 0);  -- SDRAM_Master_avalon_master_translator:uav_burstcount -> sdram_controller_s1_translator:uav_burstcount
	signal sdram_master_avalon_master_translator_avalon_universal_master_0_writedata     : std_logic_vector(31 downto 0); -- SDRAM_Master_avalon_master_translator:uav_writedata -> sdram_controller_s1_translator:uav_writedata
	signal sdram_master_avalon_master_translator_avalon_universal_master_0_address       : std_logic_vector(22 downto 0); -- SDRAM_Master_avalon_master_translator:uav_address -> sdram_controller_s1_translator:uav_address
	signal sdram_master_avalon_master_translator_avalon_universal_master_0_lock          : std_logic;                     -- SDRAM_Master_avalon_master_translator:uav_lock -> sdram_controller_s1_translator:uav_lock
	signal sdram_master_avalon_master_translator_avalon_universal_master_0_write         : std_logic;                     -- SDRAM_Master_avalon_master_translator:uav_write -> sdram_controller_s1_translator:uav_write
	signal sdram_master_avalon_master_translator_avalon_universal_master_0_read          : std_logic;                     -- SDRAM_Master_avalon_master_translator:uav_read -> sdram_controller_s1_translator:uav_read
	signal sdram_master_avalon_master_translator_avalon_universal_master_0_readdata      : std_logic_vector(31 downto 0); -- sdram_controller_s1_translator:uav_readdata -> SDRAM_Master_avalon_master_translator:uav_readdata
	signal sdram_master_avalon_master_translator_avalon_universal_master_0_debugaccess   : std_logic;                     -- SDRAM_Master_avalon_master_translator:uav_debugaccess -> sdram_controller_s1_translator:uav_debugaccess
	signal sdram_master_avalon_master_translator_avalon_universal_master_0_byteenable    : std_logic_vector(3 downto 0);  -- SDRAM_Master_avalon_master_translator:uav_byteenable -> sdram_controller_s1_translator:uav_byteenable
	signal sdram_master_avalon_master_translator_avalon_universal_master_0_readdatavalid : std_logic;                     -- sdram_controller_s1_translator:uav_readdatavalid -> SDRAM_Master_avalon_master_translator:uav_readdatavalid
	signal sdram_controller_s1_translator_avalon_anti_slave_0_waitrequest                : std_logic;                     -- sdram_controller:za_waitrequest -> sdram_controller_s1_translator:av_waitrequest
	signal sdram_controller_s1_translator_avalon_anti_slave_0_writedata                  : std_logic_vector(31 downto 0); -- sdram_controller_s1_translator:av_writedata -> sdram_controller:az_data
	signal sdram_controller_s1_translator_avalon_anti_slave_0_address                    : std_logic_vector(20 downto 0); -- sdram_controller_s1_translator:av_address -> sdram_controller:az_addr
	signal sdram_controller_s1_translator_avalon_anti_slave_0_chipselect                 : std_logic;                     -- sdram_controller_s1_translator:av_chipselect -> sdram_controller:az_cs
	signal sdram_controller_s1_translator_avalon_anti_slave_0_write                      : std_logic;                     -- sdram_controller_s1_translator:av_write -> sdram_controller_s1_translator_avalon_anti_slave_0_write:in
	signal sdram_controller_s1_translator_avalon_anti_slave_0_read                       : std_logic;                     -- sdram_controller_s1_translator:av_read -> sdram_controller_s1_translator_avalon_anti_slave_0_read:in
	signal sdram_controller_s1_translator_avalon_anti_slave_0_readdata                   : std_logic_vector(31 downto 0); -- sdram_controller:za_data -> sdram_controller_s1_translator:av_readdata
	signal sdram_controller_s1_translator_avalon_anti_slave_0_readdatavalid              : std_logic;                     -- sdram_controller:za_valid -> sdram_controller_s1_translator:av_readdatavalid
	signal sdram_controller_s1_translator_avalon_anti_slave_0_byteenable                 : std_logic_vector(3 downto 0);  -- sdram_controller_s1_translator:av_byteenable -> sdram_controller_s1_translator_avalon_anti_slave_0_byteenable:in
	signal rst_controller_reset_out_reset                                                : std_logic;                     -- rst_controller:reset_out -> [SDRAM_Master:KEY, SDRAM_Master_avalon_master_translator:reset, rst_controller_reset_out_reset:in, sdram_controller_s1_translator:reset]
	signal reset_reset_n_ports_inv                                                       : std_logic;                     -- reset_reset_n:inv -> rst_controller:reset_in0
	signal sdram_controller_s1_translator_avalon_anti_slave_0_write_ports_inv            : std_logic;                     -- sdram_controller_s1_translator_avalon_anti_slave_0_write:inv -> sdram_controller:az_wr_n
	signal sdram_controller_s1_translator_avalon_anti_slave_0_read_ports_inv             : std_logic;                     -- sdram_controller_s1_translator_avalon_anti_slave_0_read:inv -> sdram_controller:az_rd_n
	signal sdram_controller_s1_translator_avalon_anti_slave_0_byteenable_ports_inv       : std_logic_vector(3 downto 0);  -- sdram_controller_s1_translator_avalon_anti_slave_0_byteenable:inv -> sdram_controller:az_be_n
	signal rst_controller_reset_out_reset_ports_inv                                      : std_logic;                     -- rst_controller_reset_out_reset:inv -> sdram_controller:reset_n

begin

	sdram_controller : component SDRAM_sdram_controller
		port map (
			clk            => clk_clk,                                                                 --   clk.clk
			reset_n        => rst_controller_reset_out_reset_ports_inv,                                -- reset.reset_n
			az_addr        => sdram_controller_s1_translator_avalon_anti_slave_0_address,              --    s1.address
			az_be_n        => sdram_controller_s1_translator_avalon_anti_slave_0_byteenable_ports_inv, --      .byteenable_n
			az_cs          => sdram_controller_s1_translator_avalon_anti_slave_0_chipselect,           --      .chipselect
			az_data        => sdram_controller_s1_translator_avalon_anti_slave_0_writedata,            --      .writedata
			az_rd_n        => sdram_controller_s1_translator_avalon_anti_slave_0_read_ports_inv,       --      .read_n
			az_wr_n        => sdram_controller_s1_translator_avalon_anti_slave_0_write_ports_inv,      --      .write_n
			za_data        => sdram_controller_s1_translator_avalon_anti_slave_0_readdata,             --      .readdata
			za_valid       => sdram_controller_s1_translator_avalon_anti_slave_0_readdatavalid,        --      .readdatavalid
			za_waitrequest => sdram_controller_s1_translator_avalon_anti_slave_0_waitrequest,          --      .waitrequest
			zs_addr        => open,                                                                    --  wire.export
			zs_ba          => open,                                                                    --      .export
			zs_cas_n       => open,                                                                    --      .export
			zs_cke         => open,                                                                    --      .export
			zs_cs_n        => open,                                                                    --      .export
			zs_dq          => open,                                                                    --      .export
			zs_dqm         => open,                                                                    --      .export
			zs_ras_n       => open,                                                                    --      .export
			zs_we_n        => open                                                                     --      .export
		);

	sdram_master : component SDRAM_SDRAM_Master
		port map (
			CLOCK_50        => clk_clk,                                  --    clock_sink.clk
			KEY             => rst_controller_reset_out_reset,           --    reset_sink.reset
			HEX0            => open,                                     --   conduit_end.export
			HEX1            => open,                                     --              .export
			HEX3            => open,                                     --              .export
			HEX2            => open,                                     --              .export
			m_waitrequest   => sdram_master_avalon_master_waitrequest,   -- avalon_master.waitrequest
			m_readdatavalid => sdram_master_avalon_master_readdatavalid, --              .readdatavalid
			m_readdata      => sdram_master_avalon_master_readdata,      --              .readdata
			m_write         => sdram_master_avalon_master_write,         --              .write
			m_read          => sdram_master_avalon_master_read,          --              .read
			m_address       => sdram_master_avalon_master_address,       --              .address
			m_byteenable    => sdram_master_avalon_master_byteenable,    --              .byteenable
			m_writedata     => sdram_master_avalon_master_writedata      --              .writedata
		);

	sdram_master_avalon_master_translator : component altera_merlin_master_translator
		generic map (
			AV_ADDRESS_W                => 21,
			AV_DATA_W                   => 32,
			AV_BURSTCOUNT_W             => 1,
			AV_BYTEENABLE_W             => 4,
			UAV_ADDRESS_W               => 23,
			UAV_BURSTCOUNT_W            => 3,
			USE_READ                    => 1,
			USE_WRITE                   => 1,
			USE_BEGINBURSTTRANSFER      => 0,
			USE_BEGINTRANSFER           => 0,
			USE_CHIPSELECT              => 0,
			USE_BURSTCOUNT              => 0,
			USE_READDATAVALID           => 1,
			USE_WAITREQUEST             => 1,
			USE_READRESPONSE            => 0,
			USE_WRITERESPONSE           => 0,
			AV_SYMBOLS_PER_WORD         => 4,
			AV_ADDRESS_SYMBOLS          => 0,
			AV_BURSTCOUNT_SYMBOLS       => 0,
			AV_CONSTANT_BURST_BEHAVIOR  => 0,
			UAV_CONSTANT_BURST_BEHAVIOR => 0,
			AV_LINEWRAPBURSTS           => 0,
			AV_REGISTERINCOMINGSIGNALS  => 0
		)
		port map (
			clk                      => clk_clk,                                                                       --                       clk.clk
			reset                    => rst_controller_reset_out_reset,                                                --                     reset.reset
			uav_address              => sdram_master_avalon_master_translator_avalon_universal_master_0_address,       -- avalon_universal_master_0.address
			uav_burstcount           => sdram_master_avalon_master_translator_avalon_universal_master_0_burstcount,    --                          .burstcount
			uav_read                 => sdram_master_avalon_master_translator_avalon_universal_master_0_read,          --                          .read
			uav_write                => sdram_master_avalon_master_translator_avalon_universal_master_0_write,         --                          .write
			uav_waitrequest          => sdram_master_avalon_master_translator_avalon_universal_master_0_waitrequest,   --                          .waitrequest
			uav_readdatavalid        => sdram_master_avalon_master_translator_avalon_universal_master_0_readdatavalid, --                          .readdatavalid
			uav_byteenable           => sdram_master_avalon_master_translator_avalon_universal_master_0_byteenable,    --                          .byteenable
			uav_readdata             => sdram_master_avalon_master_translator_avalon_universal_master_0_readdata,      --                          .readdata
			uav_writedata            => sdram_master_avalon_master_translator_avalon_universal_master_0_writedata,     --                          .writedata
			uav_lock                 => sdram_master_avalon_master_translator_avalon_universal_master_0_lock,          --                          .lock
			uav_debugaccess          => sdram_master_avalon_master_translator_avalon_universal_master_0_debugaccess,   --                          .debugaccess
			av_address               => sdram_master_avalon_master_address,                                            --      avalon_anti_master_0.address
			av_waitrequest           => sdram_master_avalon_master_waitrequest,                                        --                          .waitrequest
			av_byteenable            => sdram_master_avalon_master_byteenable,                                         --                          .byteenable
			av_read                  => sdram_master_avalon_master_read,                                               --                          .read
			av_readdata              => sdram_master_avalon_master_readdata,                                           --                          .readdata
			av_readdatavalid         => sdram_master_avalon_master_readdatavalid,                                      --                          .readdatavalid
			av_write                 => sdram_master_avalon_master_write,                                              --                          .write
			av_writedata             => sdram_master_avalon_master_writedata,                                          --                          .writedata
			av_burstcount            => "1",                                                                           --               (terminated)
			av_beginbursttransfer    => '0',                                                                           --               (terminated)
			av_begintransfer         => '0',                                                                           --               (terminated)
			av_chipselect            => '0',                                                                           --               (terminated)
			av_lock                  => '0',                                                                           --               (terminated)
			av_debugaccess           => '0',                                                                           --               (terminated)
			uav_clken                => open,                                                                          --               (terminated)
			av_clken                 => '1',                                                                           --               (terminated)
			uav_response             => "00",                                                                          --               (terminated)
			av_response              => open,                                                                          --               (terminated)
			uav_writeresponserequest => open,                                                                          --               (terminated)
			uav_writeresponsevalid   => '0',                                                                           --               (terminated)
			av_writeresponserequest  => '0',                                                                           --               (terminated)
			av_writeresponsevalid    => open                                                                           --               (terminated)
		);

	sdram_controller_s1_translator : component altera_merlin_slave_translator
		generic map (
			AV_ADDRESS_W                   => 21,
			AV_DATA_W                      => 32,
			UAV_DATA_W                     => 32,
			AV_BURSTCOUNT_W                => 1,
			AV_BYTEENABLE_W                => 4,
			UAV_BYTEENABLE_W               => 4,
			UAV_ADDRESS_W                  => 23,
			UAV_BURSTCOUNT_W               => 3,
			AV_READLATENCY                 => 0,
			USE_READDATAVALID              => 1,
			USE_WAITREQUEST                => 1,
			USE_UAV_CLKEN                  => 0,
			USE_READRESPONSE               => 0,
			USE_WRITERESPONSE              => 0,
			AV_SYMBOLS_PER_WORD            => 4,
			AV_ADDRESS_SYMBOLS             => 0,
			AV_BURSTCOUNT_SYMBOLS          => 0,
			AV_CONSTANT_BURST_BEHAVIOR     => 0,
			UAV_CONSTANT_BURST_BEHAVIOR    => 0,
			AV_REQUIRE_UNALIGNED_ADDRESSES => 0,
			CHIPSELECT_THROUGH_READLATENCY => 0,
			AV_READ_WAIT_CYCLES            => 1,
			AV_WRITE_WAIT_CYCLES           => 0,
			AV_SETUP_WAIT_CYCLES           => 0,
			AV_DATA_HOLD_CYCLES            => 0
		)
		port map (
			clk                      => clk_clk,                                                                       --                      clk.clk
			reset                    => rst_controller_reset_out_reset,                                                --                    reset.reset
			uav_address              => sdram_master_avalon_master_translator_avalon_universal_master_0_address,       -- avalon_universal_slave_0.address
			uav_burstcount           => sdram_master_avalon_master_translator_avalon_universal_master_0_burstcount,    --                         .burstcount
			uav_read                 => sdram_master_avalon_master_translator_avalon_universal_master_0_read,          --                         .read
			uav_write                => sdram_master_avalon_master_translator_avalon_universal_master_0_write,         --                         .write
			uav_waitrequest          => sdram_master_avalon_master_translator_avalon_universal_master_0_waitrequest,   --                         .waitrequest
			uav_readdatavalid        => sdram_master_avalon_master_translator_avalon_universal_master_0_readdatavalid, --                         .readdatavalid
			uav_byteenable           => sdram_master_avalon_master_translator_avalon_universal_master_0_byteenable,    --                         .byteenable
			uav_readdata             => sdram_master_avalon_master_translator_avalon_universal_master_0_readdata,      --                         .readdata
			uav_writedata            => sdram_master_avalon_master_translator_avalon_universal_master_0_writedata,     --                         .writedata
			uav_lock                 => sdram_master_avalon_master_translator_avalon_universal_master_0_lock,          --                         .lock
			uav_debugaccess          => sdram_master_avalon_master_translator_avalon_universal_master_0_debugaccess,   --                         .debugaccess
			av_address               => sdram_controller_s1_translator_avalon_anti_slave_0_address,                    --      avalon_anti_slave_0.address
			av_write                 => sdram_controller_s1_translator_avalon_anti_slave_0_write,                      --                         .write
			av_read                  => sdram_controller_s1_translator_avalon_anti_slave_0_read,                       --                         .read
			av_readdata              => sdram_controller_s1_translator_avalon_anti_slave_0_readdata,                   --                         .readdata
			av_writedata             => sdram_controller_s1_translator_avalon_anti_slave_0_writedata,                  --                         .writedata
			av_byteenable            => sdram_controller_s1_translator_avalon_anti_slave_0_byteenable,                 --                         .byteenable
			av_readdatavalid         => sdram_controller_s1_translator_avalon_anti_slave_0_readdatavalid,              --                         .readdatavalid
			av_waitrequest           => sdram_controller_s1_translator_avalon_anti_slave_0_waitrequest,                --                         .waitrequest
			av_chipselect            => sdram_controller_s1_translator_avalon_anti_slave_0_chipselect,                 --                         .chipselect
			av_begintransfer         => open,                                                                          --              (terminated)
			av_beginbursttransfer    => open,                                                                          --              (terminated)
			av_burstcount            => open,                                                                          --              (terminated)
			av_writebyteenable       => open,                                                                          --              (terminated)
			av_lock                  => open,                                                                          --              (terminated)
			av_clken                 => open,                                                                          --              (terminated)
			uav_clken                => '0',                                                                           --              (terminated)
			av_debugaccess           => open,                                                                          --              (terminated)
			av_outputenable          => open,                                                                          --              (terminated)
			uav_response             => open,                                                                          --              (terminated)
			av_response              => "00",                                                                          --              (terminated)
			uav_writeresponserequest => '0',                                                                           --              (terminated)
			uav_writeresponsevalid   => open,                                                                          --              (terminated)
			av_writeresponserequest  => open,                                                                          --              (terminated)
			av_writeresponsevalid    => '0'                                                                            --              (terminated)
		);

	rst_controller : component altera_reset_controller
		generic map (
			NUM_RESET_INPUTS        => 1,
			OUTPUT_RESET_SYNC_EDGES => "deassert",
			SYNC_DEPTH              => 2,
			RESET_REQUEST_PRESENT   => 0
		)
		port map (
			reset_in0  => reset_reset_n_ports_inv,        -- reset_in0.reset
			clk        => clk_clk,                        --       clk.clk
			reset_out  => rst_controller_reset_out_reset, -- reset_out.reset
			reset_req  => open,                           -- (terminated)
			reset_in1  => '0',                            -- (terminated)
			reset_in2  => '0',                            -- (terminated)
			reset_in3  => '0',                            -- (terminated)
			reset_in4  => '0',                            -- (terminated)
			reset_in5  => '0',                            -- (terminated)
			reset_in6  => '0',                            -- (terminated)
			reset_in7  => '0',                            -- (terminated)
			reset_in8  => '0',                            -- (terminated)
			reset_in9  => '0',                            -- (terminated)
			reset_in10 => '0',                            -- (terminated)
			reset_in11 => '0',                            -- (terminated)
			reset_in12 => '0',                            -- (terminated)
			reset_in13 => '0',                            -- (terminated)
			reset_in14 => '0',                            -- (terminated)
			reset_in15 => '0'                             -- (terminated)
		);

	reset_reset_n_ports_inv <= not reset_reset_n;

	sdram_controller_s1_translator_avalon_anti_slave_0_write_ports_inv <= not sdram_controller_s1_translator_avalon_anti_slave_0_write;

	sdram_controller_s1_translator_avalon_anti_slave_0_read_ports_inv <= not sdram_controller_s1_translator_avalon_anti_slave_0_read;

	sdram_controller_s1_translator_avalon_anti_slave_0_byteenable_ports_inv <= not sdram_controller_s1_translator_avalon_anti_slave_0_byteenable;

	rst_controller_reset_out_reset_ports_inv <= not rst_controller_reset_out_reset;

end architecture rtl; -- of SDRAM
