-- Avalon_Blockram.vhd

-- Generated using ACDS version 13.0sp1 232 at 2016.02.05.12:16:14

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity Avalon_Blockram is
	port (
		clk_clk       : in std_logic := '0'; --   clk.clk
		reset_reset_n : in std_logic := '0'  -- reset.reset_n
	);
end entity Avalon_Blockram;

architecture rtl of Avalon_Blockram is
	component Avalon_Blockram_onchip_memory2_0 is
		port (
			clk        : in  std_logic                     := 'X';             -- clk
			address    : in  std_logic_vector(7 downto 0)  := (others => 'X'); -- address
			clken      : in  std_logic                     := 'X';             -- clken
			chipselect : in  std_logic                     := 'X';             -- chipselect
			write      : in  std_logic                     := 'X';             -- write
			readdata   : out std_logic_vector(31 downto 0);                    -- readdata
			writedata  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			byteenable : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			reset      : in  std_logic                     := 'X';             -- reset
			reset_req  : in  std_logic                     := 'X'              -- reset_req
		);
	end component Avalon_Blockram_onchip_memory2_0;

	component RISCV is
		port (
			CLOCK_50      : in  std_logic                     := 'X';             -- clk
			KEY           : in  std_logic_vector(0 downto 0)  := (others => 'X'); -- reset
			m_waitrequest : in  std_logic                     := 'X';             -- waitrequest
			m_readdata    : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			m_write       : out std_logic;                                        -- write
			m_read        : out std_logic;                                        -- read
			m_address     : out std_logic_vector(9 downto 0);                     -- address
			m_byteenable  : out std_logic_vector(3 downto 0);                     -- byteenable
			m_writedata   : out std_logic_vector(31 downto 0);                    -- writedata
			HEX0          : out std_logic_vector(6 downto 0);                     -- export
			HEX2          : out std_logic_vector(6 downto 0);                     -- export
			HEX3          : out std_logic_vector(6 downto 0);                     -- export
			HEX1          : out std_logic_vector(6 downto 0)                      -- export
		);
	end component RISCV;

	component altera_merlin_master_translator is
		generic (
			AV_ADDRESS_W                : integer := 32;
			AV_DATA_W                   : integer := 32;
			AV_BURSTCOUNT_W             : integer := 4;
			AV_BYTEENABLE_W             : integer := 4;
			UAV_ADDRESS_W               : integer := 38;
			UAV_BURSTCOUNT_W            : integer := 10;
			USE_READ                    : integer := 1;
			USE_WRITE                   : integer := 1;
			USE_BEGINBURSTTRANSFER      : integer := 0;
			USE_BEGINTRANSFER           : integer := 0;
			USE_CHIPSELECT              : integer := 0;
			USE_BURSTCOUNT              : integer := 1;
			USE_READDATAVALID           : integer := 1;
			USE_WAITREQUEST             : integer := 1;
			USE_READRESPONSE            : integer := 0;
			USE_WRITERESPONSE           : integer := 0;
			AV_SYMBOLS_PER_WORD         : integer := 4;
			AV_ADDRESS_SYMBOLS          : integer := 0;
			AV_BURSTCOUNT_SYMBOLS       : integer := 0;
			AV_CONSTANT_BURST_BEHAVIOR  : integer := 0;
			UAV_CONSTANT_BURST_BEHAVIOR : integer := 0;
			AV_LINEWRAPBURSTS           : integer := 0;
			AV_REGISTERINCOMINGSIGNALS  : integer := 0
		);
		port (
			clk                      : in  std_logic                     := 'X';             -- clk
			reset                    : in  std_logic                     := 'X';             -- reset
			uav_address              : out std_logic_vector(11 downto 0);                    -- address
			uav_burstcount           : out std_logic_vector(2 downto 0);                     -- burstcount
			uav_read                 : out std_logic;                                        -- read
			uav_write                : out std_logic;                                        -- write
			uav_waitrequest          : in  std_logic                     := 'X';             -- waitrequest
			uav_readdatavalid        : in  std_logic                     := 'X';             -- readdatavalid
			uav_byteenable           : out std_logic_vector(3 downto 0);                     -- byteenable
			uav_readdata             : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			uav_writedata            : out std_logic_vector(31 downto 0);                    -- writedata
			uav_lock                 : out std_logic;                                        -- lock
			uav_debugaccess          : out std_logic;                                        -- debugaccess
			av_address               : in  std_logic_vector(9 downto 0)  := (others => 'X'); -- address
			av_waitrequest           : out std_logic;                                        -- waitrequest
			av_byteenable            : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			av_read                  : in  std_logic                     := 'X';             -- read
			av_readdata              : out std_logic_vector(31 downto 0);                    -- readdata
			av_write                 : in  std_logic                     := 'X';             -- write
			av_writedata             : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			av_burstcount            : in  std_logic_vector(0 downto 0)  := (others => 'X'); -- burstcount
			av_beginbursttransfer    : in  std_logic                     := 'X';             -- beginbursttransfer
			av_begintransfer         : in  std_logic                     := 'X';             -- begintransfer
			av_chipselect            : in  std_logic                     := 'X';             -- chipselect
			av_readdatavalid         : out std_logic;                                        -- readdatavalid
			av_lock                  : in  std_logic                     := 'X';             -- lock
			av_debugaccess           : in  std_logic                     := 'X';             -- debugaccess
			uav_clken                : out std_logic;                                        -- clken
			av_clken                 : in  std_logic                     := 'X';             -- clken
			uav_response             : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- response
			av_response              : out std_logic_vector(1 downto 0);                     -- response
			uav_writeresponserequest : out std_logic;                                        -- writeresponserequest
			uav_writeresponsevalid   : in  std_logic                     := 'X';             -- writeresponsevalid
			av_writeresponserequest  : in  std_logic                     := 'X';             -- writeresponserequest
			av_writeresponsevalid    : out std_logic                                         -- writeresponsevalid
		);
	end component altera_merlin_master_translator;

	component altera_merlin_slave_translator is
		generic (
			AV_ADDRESS_W                   : integer := 30;
			AV_DATA_W                      : integer := 32;
			UAV_DATA_W                     : integer := 32;
			AV_BURSTCOUNT_W                : integer := 4;
			AV_BYTEENABLE_W                : integer := 4;
			UAV_BYTEENABLE_W               : integer := 4;
			UAV_ADDRESS_W                  : integer := 32;
			UAV_BURSTCOUNT_W               : integer := 4;
			AV_READLATENCY                 : integer := 0;
			USE_READDATAVALID              : integer := 1;
			USE_WAITREQUEST                : integer := 1;
			USE_UAV_CLKEN                  : integer := 0;
			USE_READRESPONSE               : integer := 0;
			USE_WRITERESPONSE              : integer := 0;
			AV_SYMBOLS_PER_WORD            : integer := 4;
			AV_ADDRESS_SYMBOLS             : integer := 0;
			AV_BURSTCOUNT_SYMBOLS          : integer := 0;
			AV_CONSTANT_BURST_BEHAVIOR     : integer := 0;
			UAV_CONSTANT_BURST_BEHAVIOR    : integer := 0;
			AV_REQUIRE_UNALIGNED_ADDRESSES : integer := 0;
			CHIPSELECT_THROUGH_READLATENCY : integer := 0;
			AV_READ_WAIT_CYCLES            : integer := 0;
			AV_WRITE_WAIT_CYCLES           : integer := 0;
			AV_SETUP_WAIT_CYCLES           : integer := 0;
			AV_DATA_HOLD_CYCLES            : integer := 0
		);
		port (
			clk                      : in  std_logic                     := 'X';             -- clk
			reset                    : in  std_logic                     := 'X';             -- reset
			uav_address              : in  std_logic_vector(11 downto 0) := (others => 'X'); -- address
			uav_burstcount           : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- burstcount
			uav_read                 : in  std_logic                     := 'X';             -- read
			uav_write                : in  std_logic                     := 'X';             -- write
			uav_waitrequest          : out std_logic;                                        -- waitrequest
			uav_readdatavalid        : out std_logic;                                        -- readdatavalid
			uav_byteenable           : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			uav_readdata             : out std_logic_vector(31 downto 0);                    -- readdata
			uav_writedata            : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			uav_lock                 : in  std_logic                     := 'X';             -- lock
			uav_debugaccess          : in  std_logic                     := 'X';             -- debugaccess
			av_address               : out std_logic_vector(7 downto 0);                     -- address
			av_write                 : out std_logic;                                        -- write
			av_readdata              : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			av_writedata             : out std_logic_vector(31 downto 0);                    -- writedata
			av_byteenable            : out std_logic_vector(3 downto 0);                     -- byteenable
			av_chipselect            : out std_logic;                                        -- chipselect
			av_clken                 : out std_logic;                                        -- clken
			av_read                  : out std_logic;                                        -- read
			av_begintransfer         : out std_logic;                                        -- begintransfer
			av_beginbursttransfer    : out std_logic;                                        -- beginbursttransfer
			av_burstcount            : out std_logic_vector(0 downto 0);                     -- burstcount
			av_readdatavalid         : in  std_logic                     := 'X';             -- readdatavalid
			av_waitrequest           : in  std_logic                     := 'X';             -- waitrequest
			av_writebyteenable       : out std_logic_vector(3 downto 0);                     -- writebyteenable
			av_lock                  : out std_logic;                                        -- lock
			uav_clken                : in  std_logic                     := 'X';             -- clken
			av_debugaccess           : out std_logic;                                        -- debugaccess
			av_outputenable          : out std_logic;                                        -- outputenable
			uav_response             : out std_logic_vector(1 downto 0);                     -- response
			av_response              : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- response
			uav_writeresponserequest : in  std_logic                     := 'X';             -- writeresponserequest
			uav_writeresponsevalid   : out std_logic;                                        -- writeresponsevalid
			av_writeresponserequest  : out std_logic;                                        -- writeresponserequest
			av_writeresponsevalid    : in  std_logic                     := 'X'              -- writeresponsevalid
		);
	end component altera_merlin_slave_translator;

	component altera_reset_controller is
		generic (
			NUM_RESET_INPUTS        : integer := 6;
			OUTPUT_RESET_SYNC_EDGES : string  := "deassert";
			SYNC_DEPTH              : integer := 2;
			RESET_REQUEST_PRESENT   : integer := 0
		);
		port (
			reset_in0  : in  std_logic := 'X'; -- reset
			clk        : in  std_logic := 'X'; -- clk
			reset_out  : out std_logic;        -- reset
			reset_req  : out std_logic;        -- reset_req
			reset_in1  : in  std_logic := 'X'; -- reset
			reset_in2  : in  std_logic := 'X'; -- reset
			reset_in3  : in  std_logic := 'X'; -- reset
			reset_in4  : in  std_logic := 'X'; -- reset
			reset_in5  : in  std_logic := 'X'; -- reset
			reset_in6  : in  std_logic := 'X'; -- reset
			reset_in7  : in  std_logic := 'X'; -- reset
			reset_in8  : in  std_logic := 'X'; -- reset
			reset_in9  : in  std_logic := 'X'; -- reset
			reset_in10 : in  std_logic := 'X'; -- reset
			reset_in11 : in  std_logic := 'X'; -- reset
			reset_in12 : in  std_logic := 'X'; -- reset
			reset_in13 : in  std_logic := 'X'; -- reset
			reset_in14 : in  std_logic := 'X'; -- reset
			reset_in15 : in  std_logic := 'X'  -- reset
		);
	end component altera_reset_controller;

	signal blockram_masterinterface_0_avalon_master_waitrequest                                        : std_logic;                     -- Blockram_MasterInterface_0_avalon_master_translator:av_waitrequest -> Blockram_MasterInterface_0:m_waitrequest
	signal blockram_masterinterface_0_avalon_master_writedata                                          : std_logic_vector(31 downto 0); -- Blockram_MasterInterface_0:m_writedata -> Blockram_MasterInterface_0_avalon_master_translator:av_writedata
	signal blockram_masterinterface_0_avalon_master_address                                            : std_logic_vector(9 downto 0);  -- Blockram_MasterInterface_0:m_address -> Blockram_MasterInterface_0_avalon_master_translator:av_address
	signal blockram_masterinterface_0_avalon_master_write                                              : std_logic;                     -- Blockram_MasterInterface_0:m_write -> Blockram_MasterInterface_0_avalon_master_translator:av_write
	signal blockram_masterinterface_0_avalon_master_read                                               : std_logic;                     -- Blockram_MasterInterface_0:m_read -> Blockram_MasterInterface_0_avalon_master_translator:av_read
	signal blockram_masterinterface_0_avalon_master_readdata                                           : std_logic_vector(31 downto 0); -- Blockram_MasterInterface_0_avalon_master_translator:av_readdata -> Blockram_MasterInterface_0:m_readdata
	signal blockram_masterinterface_0_avalon_master_byteenable                                         : std_logic_vector(3 downto 0);  -- Blockram_MasterInterface_0:m_byteenable -> Blockram_MasterInterface_0_avalon_master_translator:av_byteenable
	signal blockram_masterinterface_0_avalon_master_translator_avalon_universal_master_0_waitrequest   : std_logic;                     -- onchip_memory2_0_s1_translator:uav_waitrequest -> Blockram_MasterInterface_0_avalon_master_translator:uav_waitrequest
	signal blockram_masterinterface_0_avalon_master_translator_avalon_universal_master_0_burstcount    : std_logic_vector(2 downto 0);  -- Blockram_MasterInterface_0_avalon_master_translator:uav_burstcount -> onchip_memory2_0_s1_translator:uav_burstcount
	signal blockram_masterinterface_0_avalon_master_translator_avalon_universal_master_0_writedata     : std_logic_vector(31 downto 0); -- Blockram_MasterInterface_0_avalon_master_translator:uav_writedata -> onchip_memory2_0_s1_translator:uav_writedata
	signal blockram_masterinterface_0_avalon_master_translator_avalon_universal_master_0_address       : std_logic_vector(11 downto 0); -- Blockram_MasterInterface_0_avalon_master_translator:uav_address -> onchip_memory2_0_s1_translator:uav_address
	signal blockram_masterinterface_0_avalon_master_translator_avalon_universal_master_0_lock          : std_logic;                     -- Blockram_MasterInterface_0_avalon_master_translator:uav_lock -> onchip_memory2_0_s1_translator:uav_lock
	signal blockram_masterinterface_0_avalon_master_translator_avalon_universal_master_0_write         : std_logic;                     -- Blockram_MasterInterface_0_avalon_master_translator:uav_write -> onchip_memory2_0_s1_translator:uav_write
	signal blockram_masterinterface_0_avalon_master_translator_avalon_universal_master_0_read          : std_logic;                     -- Blockram_MasterInterface_0_avalon_master_translator:uav_read -> onchip_memory2_0_s1_translator:uav_read
	signal blockram_masterinterface_0_avalon_master_translator_avalon_universal_master_0_readdata      : std_logic_vector(31 downto 0); -- onchip_memory2_0_s1_translator:uav_readdata -> Blockram_MasterInterface_0_avalon_master_translator:uav_readdata
	signal blockram_masterinterface_0_avalon_master_translator_avalon_universal_master_0_debugaccess   : std_logic;                     -- Blockram_MasterInterface_0_avalon_master_translator:uav_debugaccess -> onchip_memory2_0_s1_translator:uav_debugaccess
	signal blockram_masterinterface_0_avalon_master_translator_avalon_universal_master_0_byteenable    : std_logic_vector(3 downto 0);  -- Blockram_MasterInterface_0_avalon_master_translator:uav_byteenable -> onchip_memory2_0_s1_translator:uav_byteenable
	signal blockram_masterinterface_0_avalon_master_translator_avalon_universal_master_0_readdatavalid : std_logic;                     -- onchip_memory2_0_s1_translator:uav_readdatavalid -> Blockram_MasterInterface_0_avalon_master_translator:uav_readdatavalid
	signal onchip_memory2_0_s1_translator_avalon_anti_slave_0_writedata                                : std_logic_vector(31 downto 0); -- onchip_memory2_0_s1_translator:av_writedata -> onchip_memory2_0:writedata
	signal onchip_memory2_0_s1_translator_avalon_anti_slave_0_address                                  : std_logic_vector(7 downto 0);  -- onchip_memory2_0_s1_translator:av_address -> onchip_memory2_0:address
	signal onchip_memory2_0_s1_translator_avalon_anti_slave_0_chipselect                               : std_logic;                     -- onchip_memory2_0_s1_translator:av_chipselect -> onchip_memory2_0:chipselect
	signal onchip_memory2_0_s1_translator_avalon_anti_slave_0_clken                                    : std_logic;                     -- onchip_memory2_0_s1_translator:av_clken -> onchip_memory2_0:clken
	signal onchip_memory2_0_s1_translator_avalon_anti_slave_0_write                                    : std_logic;                     -- onchip_memory2_0_s1_translator:av_write -> onchip_memory2_0:write
	signal onchip_memory2_0_s1_translator_avalon_anti_slave_0_readdata                                 : std_logic_vector(31 downto 0); -- onchip_memory2_0:readdata -> onchip_memory2_0_s1_translator:av_readdata
	signal onchip_memory2_0_s1_translator_avalon_anti_slave_0_byteenable                               : std_logic_vector(3 downto 0);  -- onchip_memory2_0_s1_translator:av_byteenable -> onchip_memory2_0:byteenable
	signal rst_controller_reset_out_reset                                                              : std_logic;                     -- rst_controller:reset_out -> [Blockram_MasterInterface_0:KEY, Blockram_MasterInterface_0_avalon_master_translator:reset, onchip_memory2_0:reset, onchip_memory2_0_s1_translator:reset]
	signal rst_controller_reset_out_reset_req                                                          : std_logic;                     -- rst_controller:reset_req -> onchip_memory2_0:reset_req
	signal reset_reset_n_ports_inv                                                                     : std_logic;                     -- reset_reset_n:inv -> rst_controller:reset_in0

begin

	onchip_memory2_0 : component Avalon_Blockram_onchip_memory2_0
		port map (
			clk        => clk_clk,                                                       --   clk1.clk
			address    => onchip_memory2_0_s1_translator_avalon_anti_slave_0_address,    --     s1.address
			clken      => onchip_memory2_0_s1_translator_avalon_anti_slave_0_clken,      --       .clken
			chipselect => onchip_memory2_0_s1_translator_avalon_anti_slave_0_chipselect, --       .chipselect
			write      => onchip_memory2_0_s1_translator_avalon_anti_slave_0_write,      --       .write
			readdata   => onchip_memory2_0_s1_translator_avalon_anti_slave_0_readdata,   --       .readdata
			writedata  => onchip_memory2_0_s1_translator_avalon_anti_slave_0_writedata,  --       .writedata
			byteenable => onchip_memory2_0_s1_translator_avalon_anti_slave_0_byteenable, --       .byteenable
			reset      => rst_controller_reset_out_reset,                                -- reset1.reset
			reset_req  => rst_controller_reset_out_reset_req                             --       .reset_req
		);

	blockram_masterinterface_0 : component RISCV
		port map (
			CLOCK_50      => clk_clk,                                              --    clock_sink.clk
			KEY(0)        => rst_controller_reset_out_reset,                       --    reset_sink.reset
			m_waitrequest => blockram_masterinterface_0_avalon_master_waitrequest, -- avalon_master.waitrequest
			m_readdata    => blockram_masterinterface_0_avalon_master_readdata,    --              .readdata
			m_write       => blockram_masterinterface_0_avalon_master_write,       --              .write
			m_read        => blockram_masterinterface_0_avalon_master_read,        --              .read
			m_address     => blockram_masterinterface_0_avalon_master_address,     --              .address
			m_byteenable  => blockram_masterinterface_0_avalon_master_byteenable,  --              .byteenable
			m_writedata   => blockram_masterinterface_0_avalon_master_writedata,   --              .writedata
			HEX0          => open,                                                 --   conduit_end.export
			HEX2          => open,                                                 --              .export
			HEX3          => open,                                                 --              .export
			HEX1          => open                                                  --              .export
		);

	blockram_masterinterface_0_avalon_master_translator : component altera_merlin_master_translator
		generic map (
			AV_ADDRESS_W                => 10,
			AV_DATA_W                   => 32,
			AV_BURSTCOUNT_W             => 1,
			AV_BYTEENABLE_W             => 4,
			UAV_ADDRESS_W               => 12,
			UAV_BURSTCOUNT_W            => 3,
			USE_READ                    => 1,
			USE_WRITE                   => 1,
			USE_BEGINBURSTTRANSFER      => 0,
			USE_BEGINTRANSFER           => 0,
			USE_CHIPSELECT              => 0,
			USE_BURSTCOUNT              => 0,
			USE_READDATAVALID           => 0,
			USE_WAITREQUEST             => 1,
			USE_READRESPONSE            => 0,
			USE_WRITERESPONSE           => 0,
			AV_SYMBOLS_PER_WORD         => 4,
			AV_ADDRESS_SYMBOLS          => 0,
			AV_BURSTCOUNT_SYMBOLS       => 0,
			AV_CONSTANT_BURST_BEHAVIOR  => 0,
			UAV_CONSTANT_BURST_BEHAVIOR => 0,
			AV_LINEWRAPBURSTS           => 0,
			AV_REGISTERINCOMINGSIGNALS  => 0
		)
		port map (
			clk                      => clk_clk,                                                                                     --                       clk.clk
			reset                    => rst_controller_reset_out_reset,                                                              --                     reset.reset
			uav_address              => blockram_masterinterface_0_avalon_master_translator_avalon_universal_master_0_address,       -- avalon_universal_master_0.address
			uav_burstcount           => blockram_masterinterface_0_avalon_master_translator_avalon_universal_master_0_burstcount,    --                          .burstcount
			uav_read                 => blockram_masterinterface_0_avalon_master_translator_avalon_universal_master_0_read,          --                          .read
			uav_write                => blockram_masterinterface_0_avalon_master_translator_avalon_universal_master_0_write,         --                          .write
			uav_waitrequest          => blockram_masterinterface_0_avalon_master_translator_avalon_universal_master_0_waitrequest,   --                          .waitrequest
			uav_readdatavalid        => blockram_masterinterface_0_avalon_master_translator_avalon_universal_master_0_readdatavalid, --                          .readdatavalid
			uav_byteenable           => blockram_masterinterface_0_avalon_master_translator_avalon_universal_master_0_byteenable,    --                          .byteenable
			uav_readdata             => blockram_masterinterface_0_avalon_master_translator_avalon_universal_master_0_readdata,      --                          .readdata
			uav_writedata            => blockram_masterinterface_0_avalon_master_translator_avalon_universal_master_0_writedata,     --                          .writedata
			uav_lock                 => blockram_masterinterface_0_avalon_master_translator_avalon_universal_master_0_lock,          --                          .lock
			uav_debugaccess          => blockram_masterinterface_0_avalon_master_translator_avalon_universal_master_0_debugaccess,   --                          .debugaccess
			av_address               => blockram_masterinterface_0_avalon_master_address,                                            --      avalon_anti_master_0.address
			av_waitrequest           => blockram_masterinterface_0_avalon_master_waitrequest,                                        --                          .waitrequest
			av_byteenable            => blockram_masterinterface_0_avalon_master_byteenable,                                         --                          .byteenable
			av_read                  => blockram_masterinterface_0_avalon_master_read,                                               --                          .read
			av_readdata              => blockram_masterinterface_0_avalon_master_readdata,                                           --                          .readdata
			av_write                 => blockram_masterinterface_0_avalon_master_write,                                              --                          .write
			av_writedata             => blockram_masterinterface_0_avalon_master_writedata,                                          --                          .writedata
			av_burstcount            => "1",                                                                                         --               (terminated)
			av_beginbursttransfer    => '0',                                                                                         --               (terminated)
			av_begintransfer         => '0',                                                                                         --               (terminated)
			av_chipselect            => '0',                                                                                         --               (terminated)
			av_readdatavalid         => open,                                                                                        --               (terminated)
			av_lock                  => '0',                                                                                         --               (terminated)
			av_debugaccess           => '0',                                                                                         --               (terminated)
			uav_clken                => open,                                                                                        --               (terminated)
			av_clken                 => '1',                                                                                         --               (terminated)
			uav_response             => "00",                                                                                        --               (terminated)
			av_response              => open,                                                                                        --               (terminated)
			uav_writeresponserequest => open,                                                                                        --               (terminated)
			uav_writeresponsevalid   => '0',                                                                                         --               (terminated)
			av_writeresponserequest  => '0',                                                                                         --               (terminated)
			av_writeresponsevalid    => open                                                                                         --               (terminated)
		);

	onchip_memory2_0_s1_translator : component altera_merlin_slave_translator
		generic map (
			AV_ADDRESS_W                   => 8,
			AV_DATA_W                      => 32,
			UAV_DATA_W                     => 32,
			AV_BURSTCOUNT_W                => 1,
			AV_BYTEENABLE_W                => 4,
			UAV_BYTEENABLE_W               => 4,
			UAV_ADDRESS_W                  => 12,
			UAV_BURSTCOUNT_W               => 3,
			AV_READLATENCY                 => 1,
			USE_READDATAVALID              => 0,
			USE_WAITREQUEST                => 0,
			USE_UAV_CLKEN                  => 0,
			USE_READRESPONSE               => 0,
			USE_WRITERESPONSE              => 0,
			AV_SYMBOLS_PER_WORD            => 4,
			AV_ADDRESS_SYMBOLS             => 0,
			AV_BURSTCOUNT_SYMBOLS          => 0,
			AV_CONSTANT_BURST_BEHAVIOR     => 0,
			UAV_CONSTANT_BURST_BEHAVIOR    => 0,
			AV_REQUIRE_UNALIGNED_ADDRESSES => 0,
			CHIPSELECT_THROUGH_READLATENCY => 0,
			AV_READ_WAIT_CYCLES            => 0,
			AV_WRITE_WAIT_CYCLES           => 0,
			AV_SETUP_WAIT_CYCLES           => 0,
			AV_DATA_HOLD_CYCLES            => 0
		)
		port map (
			clk                      => clk_clk,                                                                                     --                      clk.clk
			reset                    => rst_controller_reset_out_reset,                                                              --                    reset.reset
			uav_address              => blockram_masterinterface_0_avalon_master_translator_avalon_universal_master_0_address,       -- avalon_universal_slave_0.address
			uav_burstcount           => blockram_masterinterface_0_avalon_master_translator_avalon_universal_master_0_burstcount,    --                         .burstcount
			uav_read                 => blockram_masterinterface_0_avalon_master_translator_avalon_universal_master_0_read,          --                         .read
			uav_write                => blockram_masterinterface_0_avalon_master_translator_avalon_universal_master_0_write,         --                         .write
			uav_waitrequest          => blockram_masterinterface_0_avalon_master_translator_avalon_universal_master_0_waitrequest,   --                         .waitrequest
			uav_readdatavalid        => blockram_masterinterface_0_avalon_master_translator_avalon_universal_master_0_readdatavalid, --                         .readdatavalid
			uav_byteenable           => blockram_masterinterface_0_avalon_master_translator_avalon_universal_master_0_byteenable,    --                         .byteenable
			uav_readdata             => blockram_masterinterface_0_avalon_master_translator_avalon_universal_master_0_readdata,      --                         .readdata
			uav_writedata            => blockram_masterinterface_0_avalon_master_translator_avalon_universal_master_0_writedata,     --                         .writedata
			uav_lock                 => blockram_masterinterface_0_avalon_master_translator_avalon_universal_master_0_lock,          --                         .lock
			uav_debugaccess          => blockram_masterinterface_0_avalon_master_translator_avalon_universal_master_0_debugaccess,   --                         .debugaccess
			av_address               => onchip_memory2_0_s1_translator_avalon_anti_slave_0_address,                                  --      avalon_anti_slave_0.address
			av_write                 => onchip_memory2_0_s1_translator_avalon_anti_slave_0_write,                                    --                         .write
			av_readdata              => onchip_memory2_0_s1_translator_avalon_anti_slave_0_readdata,                                 --                         .readdata
			av_writedata             => onchip_memory2_0_s1_translator_avalon_anti_slave_0_writedata,                                --                         .writedata
			av_byteenable            => onchip_memory2_0_s1_translator_avalon_anti_slave_0_byteenable,                               --                         .byteenable
			av_chipselect            => onchip_memory2_0_s1_translator_avalon_anti_slave_0_chipselect,                               --                         .chipselect
			av_clken                 => onchip_memory2_0_s1_translator_avalon_anti_slave_0_clken,                                    --                         .clken
			av_read                  => open,                                                                                        --              (terminated)
			av_begintransfer         => open,                                                                                        --              (terminated)
			av_beginbursttransfer    => open,                                                                                        --              (terminated)
			av_burstcount            => open,                                                                                        --              (terminated)
			av_readdatavalid         => '0',                                                                                         --              (terminated)
			av_waitrequest           => '0',                                                                                         --              (terminated)
			av_writebyteenable       => open,                                                                                        --              (terminated)
			av_lock                  => open,                                                                                        --              (terminated)
			uav_clken                => '0',                                                                                         --              (terminated)
			av_debugaccess           => open,                                                                                        --              (terminated)
			av_outputenable          => open,                                                                                        --              (terminated)
			uav_response             => open,                                                                                        --              (terminated)
			av_response              => "00",                                                                                        --              (terminated)
			uav_writeresponserequest => '0',                                                                                         --              (terminated)
			uav_writeresponsevalid   => open,                                                                                        --              (terminated)
			av_writeresponserequest  => open,                                                                                        --              (terminated)
			av_writeresponsevalid    => '0'                                                                                          --              (terminated)
		);

	rst_controller : component altera_reset_controller
		generic map (
			NUM_RESET_INPUTS        => 1,
			OUTPUT_RESET_SYNC_EDGES => "deassert",
			SYNC_DEPTH              => 2,
			RESET_REQUEST_PRESENT   => 1
		)
		port map (
			reset_in0  => reset_reset_n_ports_inv,            -- reset_in0.reset
			clk        => clk_clk,                            --       clk.clk
			reset_out  => rst_controller_reset_out_reset,     -- reset_out.reset
			reset_req  => rst_controller_reset_out_reset_req, --          .reset_req
			reset_in1  => '0',                                -- (terminated)
			reset_in2  => '0',                                -- (terminated)
			reset_in3  => '0',                                -- (terminated)
			reset_in4  => '0',                                -- (terminated)
			reset_in5  => '0',                                -- (terminated)
			reset_in6  => '0',                                -- (terminated)
			reset_in7  => '0',                                -- (terminated)
			reset_in8  => '0',                                -- (terminated)
			reset_in9  => '0',                                -- (terminated)
			reset_in10 => '0',                                -- (terminated)
			reset_in11 => '0',                                -- (terminated)
			reset_in12 => '0',                                -- (terminated)
			reset_in13 => '0',                                -- (terminated)
			reset_in14 => '0',                                -- (terminated)
			reset_in15 => '0'                                 -- (terminated)
		);

	reset_reset_n_ports_inv <= not reset_reset_n;

end architecture rtl; -- of Avalon_Blockram
