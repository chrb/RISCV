-- FetchMemory_Blockram.vhd

-- Generated using ACDS version 13.0sp1 232 at 2016.02.03.18:27:34

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity FetchMemory_Blockram is
	port (
		clk_clk       : in std_logic := '0'; --   clk.clk
		reset_reset_n : in std_logic := '0'  -- reset.reset_n
	);
end entity FetchMemory_Blockram;

architecture rtl of FetchMemory_Blockram is
	component FetchMemory_Blockram_Memory is
		port (
			clk        : in  std_logic                     := 'X';             -- clk
			address    : in  std_logic_vector(9 downto 0)  := (others => 'X'); -- address
			clken      : in  std_logic                     := 'X';             -- clken
			chipselect : in  std_logic                     := 'X';             -- chipselect
			write      : in  std_logic                     := 'X';             -- write
			readdata   : out std_logic_vector(31 downto 0);                    -- readdata
			writedata  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			byteenable : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			reset      : in  std_logic                     := 'X';             -- reset
			reset_req  : in  std_logic                     := 'X'              -- reset_req
		);
	end component FetchMemory_Blockram_Memory;

	component FetchMemory_Blockram_InstructionMemory is
		port (
			clk         : in  std_logic                     := 'X';             -- clk
			address     : in  std_logic_vector(9 downto 0)  := (others => 'X'); -- address
			debugaccess : in  std_logic                     := 'X';             -- debugaccess
			clken       : in  std_logic                     := 'X';             -- clken
			chipselect  : in  std_logic                     := 'X';             -- chipselect
			write       : in  std_logic                     := 'X';             -- write
			readdata    : out std_logic_vector(31 downto 0);                    -- readdata
			writedata   : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			byteenable  : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			reset       : in  std_logic                     := 'X';             -- reset
			reset_req   : in  std_logic                     := 'X'              -- reset_req
		);
	end component FetchMemory_Blockram_InstructionMemory;

	component RISCV is
		port (
			CLOCK_50          : in  std_logic                     := 'X';             -- clk
			KEY               : in  std_logic_vector(0 downto 0)  := (others => 'X'); -- reset
			fetch_waitrequest : in  std_logic                     := 'X';             -- waitrequest
			fetch_readdata    : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			fetch_read        : out std_logic;                                        -- read
			fetch_address     : out std_logic_vector(9 downto 0);                     -- address
			fetch_byteenable  : out std_logic_vector(3 downto 0);                     -- byteenable
			m_waitrequest     : in  std_logic                     := 'X';             -- waitrequest
			m_readdata        : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			m_write           : out std_logic;                                        -- write
			m_read            : out std_logic;                                        -- read
			m_address         : out std_logic_vector(9 downto 0);                     -- address
			m_byteenable      : out std_logic_vector(3 downto 0);                     -- byteenable
			m_writedata       : out std_logic_vector(31 downto 0);                    -- writedata
			HEX0              : out std_logic_vector(6 downto 0);                     -- export
			HEX1              : out std_logic_vector(6 downto 0);                     -- export
			HEX2              : out std_logic_vector(6 downto 0);                     -- export
			HEX3              : out std_logic_vector(6 downto 0)                      -- export
		);
	end component RISCV;

	component fetchmemory_blockram_instructionmemory_s1_translator is
		generic (
			AV_ADDRESS_W                   : integer := 30;
			AV_DATA_W                      : integer := 32;
			UAV_DATA_W                     : integer := 32;
			AV_BURSTCOUNT_W                : integer := 4;
			AV_BYTEENABLE_W                : integer := 4;
			UAV_BYTEENABLE_W               : integer := 4;
			UAV_ADDRESS_W                  : integer := 32;
			UAV_BURSTCOUNT_W               : integer := 4;
			AV_READLATENCY                 : integer := 0;
			USE_READDATAVALID              : integer := 1;
			USE_WAITREQUEST                : integer := 1;
			USE_UAV_CLKEN                  : integer := 0;
			USE_READRESPONSE               : integer := 0;
			USE_WRITERESPONSE              : integer := 0;
			AV_SYMBOLS_PER_WORD            : integer := 4;
			AV_ADDRESS_SYMBOLS             : integer := 0;
			AV_BURSTCOUNT_SYMBOLS          : integer := 0;
			AV_CONSTANT_BURST_BEHAVIOR     : integer := 0;
			UAV_CONSTANT_BURST_BEHAVIOR    : integer := 0;
			AV_REQUIRE_UNALIGNED_ADDRESSES : integer := 0;
			CHIPSELECT_THROUGH_READLATENCY : integer := 0;
			AV_READ_WAIT_CYCLES            : integer := 0;
			AV_WRITE_WAIT_CYCLES           : integer := 0;
			AV_SETUP_WAIT_CYCLES           : integer := 0;
			AV_DATA_HOLD_CYCLES            : integer := 0
		);
		port (
			clk                      : in  std_logic                     := 'X';             -- clk
			reset                    : in  std_logic                     := 'X';             -- reset
			uav_address              : in  std_logic_vector(11 downto 0) := (others => 'X'); -- address
			uav_burstcount           : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- burstcount
			uav_read                 : in  std_logic                     := 'X';             -- read
			uav_write                : in  std_logic                     := 'X';             -- write
			uav_waitrequest          : out std_logic;                                        -- waitrequest
			uav_readdatavalid        : out std_logic;                                        -- readdatavalid
			uav_byteenable           : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			uav_readdata             : out std_logic_vector(31 downto 0);                    -- readdata
			uav_writedata            : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			uav_lock                 : in  std_logic                     := 'X';             -- lock
			uav_debugaccess          : in  std_logic                     := 'X';             -- debugaccess
			av_address               : out std_logic_vector(9 downto 0);                     -- address
			av_write                 : out std_logic;                                        -- write
			av_readdata              : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			av_writedata             : out std_logic_vector(31 downto 0);                    -- writedata
			av_byteenable            : out std_logic_vector(3 downto 0);                     -- byteenable
			av_chipselect            : out std_logic;                                        -- chipselect
			av_clken                 : out std_logic;                                        -- clken
			av_debugaccess           : out std_logic;                                        -- debugaccess
			av_read                  : out std_logic;                                        -- read
			av_begintransfer         : out std_logic;                                        -- begintransfer
			av_beginbursttransfer    : out std_logic;                                        -- beginbursttransfer
			av_burstcount            : out std_logic_vector(0 downto 0);                     -- burstcount
			av_readdatavalid         : in  std_logic                     := 'X';             -- readdatavalid
			av_waitrequest           : in  std_logic                     := 'X';             -- waitrequest
			av_writebyteenable       : out std_logic_vector(3 downto 0);                     -- writebyteenable
			av_lock                  : out std_logic;                                        -- lock
			uav_clken                : in  std_logic                     := 'X';             -- clken
			av_outputenable          : out std_logic;                                        -- outputenable
			uav_response             : out std_logic_vector(1 downto 0);                     -- response
			av_response              : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- response
			uav_writeresponserequest : in  std_logic                     := 'X';             -- writeresponserequest
			uav_writeresponsevalid   : out std_logic;                                        -- writeresponsevalid
			av_writeresponserequest  : out std_logic;                                        -- writeresponserequest
			av_writeresponsevalid    : in  std_logic                     := 'X'              -- writeresponsevalid
		);
	end component fetchmemory_blockram_instructionmemory_s1_translator;

	component fetchmemory_blockram_memory_s1_translator is
		generic (
			AV_ADDRESS_W                   : integer := 30;
			AV_DATA_W                      : integer := 32;
			UAV_DATA_W                     : integer := 32;
			AV_BURSTCOUNT_W                : integer := 4;
			AV_BYTEENABLE_W                : integer := 4;
			UAV_BYTEENABLE_W               : integer := 4;
			UAV_ADDRESS_W                  : integer := 32;
			UAV_BURSTCOUNT_W               : integer := 4;
			AV_READLATENCY                 : integer := 0;
			USE_READDATAVALID              : integer := 1;
			USE_WAITREQUEST                : integer := 1;
			USE_UAV_CLKEN                  : integer := 0;
			USE_READRESPONSE               : integer := 0;
			USE_WRITERESPONSE              : integer := 0;
			AV_SYMBOLS_PER_WORD            : integer := 4;
			AV_ADDRESS_SYMBOLS             : integer := 0;
			AV_BURSTCOUNT_SYMBOLS          : integer := 0;
			AV_CONSTANT_BURST_BEHAVIOR     : integer := 0;
			UAV_CONSTANT_BURST_BEHAVIOR    : integer := 0;
			AV_REQUIRE_UNALIGNED_ADDRESSES : integer := 0;
			CHIPSELECT_THROUGH_READLATENCY : integer := 0;
			AV_READ_WAIT_CYCLES            : integer := 0;
			AV_WRITE_WAIT_CYCLES           : integer := 0;
			AV_SETUP_WAIT_CYCLES           : integer := 0;
			AV_DATA_HOLD_CYCLES            : integer := 0
		);
		port (
			clk                      : in  std_logic                     := 'X';             -- clk
			reset                    : in  std_logic                     := 'X';             -- reset
			uav_address              : in  std_logic_vector(11 downto 0) := (others => 'X'); -- address
			uav_burstcount           : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- burstcount
			uav_read                 : in  std_logic                     := 'X';             -- read
			uav_write                : in  std_logic                     := 'X';             -- write
			uav_waitrequest          : out std_logic;                                        -- waitrequest
			uav_readdatavalid        : out std_logic;                                        -- readdatavalid
			uav_byteenable           : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			uav_readdata             : out std_logic_vector(31 downto 0);                    -- readdata
			uav_writedata            : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			uav_lock                 : in  std_logic                     := 'X';             -- lock
			uav_debugaccess          : in  std_logic                     := 'X';             -- debugaccess
			av_address               : out std_logic_vector(9 downto 0);                     -- address
			av_write                 : out std_logic;                                        -- write
			av_readdata              : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			av_writedata             : out std_logic_vector(31 downto 0);                    -- writedata
			av_byteenable            : out std_logic_vector(3 downto 0);                     -- byteenable
			av_chipselect            : out std_logic;                                        -- chipselect
			av_clken                 : out std_logic;                                        -- clken
			av_read                  : out std_logic;                                        -- read
			av_begintransfer         : out std_logic;                                        -- begintransfer
			av_beginbursttransfer    : out std_logic;                                        -- beginbursttransfer
			av_burstcount            : out std_logic_vector(0 downto 0);                     -- burstcount
			av_readdatavalid         : in  std_logic                     := 'X';             -- readdatavalid
			av_waitrequest           : in  std_logic                     := 'X';             -- waitrequest
			av_writebyteenable       : out std_logic_vector(3 downto 0);                     -- writebyteenable
			av_lock                  : out std_logic;                                        -- lock
			uav_clken                : in  std_logic                     := 'X';             -- clken
			av_debugaccess           : out std_logic;                                        -- debugaccess
			av_outputenable          : out std_logic;                                        -- outputenable
			uav_response             : out std_logic_vector(1 downto 0);                     -- response
			av_response              : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- response
			uav_writeresponserequest : in  std_logic                     := 'X';             -- writeresponserequest
			uav_writeresponsevalid   : out std_logic;                                        -- writeresponsevalid
			av_writeresponserequest  : out std_logic;                                        -- writeresponserequest
			av_writeresponsevalid    : in  std_logic                     := 'X'              -- writeresponsevalid
		);
	end component fetchmemory_blockram_memory_s1_translator;

	component fetchmemory_blockram_rst_controller is
		generic (
			NUM_RESET_INPUTS        : integer := 6;
			OUTPUT_RESET_SYNC_EDGES : string  := "deassert";
			SYNC_DEPTH              : integer := 2;
			RESET_REQUEST_PRESENT   : integer := 0
		);
		port (
			reset_in0  : in  std_logic := 'X'; -- reset
			clk        : in  std_logic := 'X'; -- clk
			reset_out  : out std_logic;        -- reset
			reset_req  : out std_logic;        -- reset_req
			reset_in1  : in  std_logic := 'X'; -- reset
			reset_in2  : in  std_logic := 'X'; -- reset
			reset_in3  : in  std_logic := 'X'; -- reset
			reset_in4  : in  std_logic := 'X'; -- reset
			reset_in5  : in  std_logic := 'X'; -- reset
			reset_in6  : in  std_logic := 'X'; -- reset
			reset_in7  : in  std_logic := 'X'; -- reset
			reset_in8  : in  std_logic := 'X'; -- reset
			reset_in9  : in  std_logic := 'X'; -- reset
			reset_in10 : in  std_logic := 'X'; -- reset
			reset_in11 : in  std_logic := 'X'; -- reset
			reset_in12 : in  std_logic := 'X'; -- reset
			reset_in13 : in  std_logic := 'X'; -- reset
			reset_in14 : in  std_logic := 'X'; -- reset
			reset_in15 : in  std_logic := 'X'  -- reset
		);
	end component fetchmemory_blockram_rst_controller;

	component fetchmemory_blockram_rst_controller_001 is
		generic (
			NUM_RESET_INPUTS        : integer := 6;
			OUTPUT_RESET_SYNC_EDGES : string  := "deassert";
			SYNC_DEPTH              : integer := 2;
			RESET_REQUEST_PRESENT   : integer := 0
		);
		port (
			reset_in0  : in  std_logic := 'X'; -- reset
			clk        : in  std_logic := 'X'; -- clk
			reset_out  : out std_logic;        -- reset
			reset_req  : out std_logic;        -- reset_req
			reset_in1  : in  std_logic := 'X'; -- reset
			reset_in2  : in  std_logic := 'X'; -- reset
			reset_in3  : in  std_logic := 'X'; -- reset
			reset_in4  : in  std_logic := 'X'; -- reset
			reset_in5  : in  std_logic := 'X'; -- reset
			reset_in6  : in  std_logic := 'X'; -- reset
			reset_in7  : in  std_logic := 'X'; -- reset
			reset_in8  : in  std_logic := 'X'; -- reset
			reset_in9  : in  std_logic := 'X'; -- reset
			reset_in10 : in  std_logic := 'X'; -- reset
			reset_in11 : in  std_logic := 'X'; -- reset
			reset_in12 : in  std_logic := 'X'; -- reset
			reset_in13 : in  std_logic := 'X'; -- reset
			reset_in14 : in  std_logic := 'X'; -- reset
			reset_in15 : in  std_logic := 'X'  -- reset
		);
	end component fetchmemory_blockram_rst_controller_001;

	component fetchmemory_blockram_masterinterface_0_fetchmaster_translator is
		generic (
			AV_ADDRESS_W                : integer := 32;
			AV_DATA_W                   : integer := 32;
			AV_BURSTCOUNT_W             : integer := 4;
			AV_BYTEENABLE_W             : integer := 4;
			UAV_ADDRESS_W               : integer := 38;
			UAV_BURSTCOUNT_W            : integer := 10;
			USE_READ                    : integer := 1;
			USE_WRITE                   : integer := 1;
			USE_BEGINBURSTTRANSFER      : integer := 0;
			USE_BEGINTRANSFER           : integer := 0;
			USE_CHIPSELECT              : integer := 0;
			USE_BURSTCOUNT              : integer := 1;
			USE_READDATAVALID           : integer := 1;
			USE_WAITREQUEST             : integer := 1;
			USE_READRESPONSE            : integer := 0;
			USE_WRITERESPONSE           : integer := 0;
			AV_SYMBOLS_PER_WORD         : integer := 4;
			AV_ADDRESS_SYMBOLS          : integer := 0;
			AV_BURSTCOUNT_SYMBOLS       : integer := 0;
			AV_CONSTANT_BURST_BEHAVIOR  : integer := 0;
			UAV_CONSTANT_BURST_BEHAVIOR : integer := 0;
			AV_LINEWRAPBURSTS           : integer := 0;
			AV_REGISTERINCOMINGSIGNALS  : integer := 0
		);
		port (
			clk                      : in  std_logic                     := 'X';             -- clk
			reset                    : in  std_logic                     := 'X';             -- reset
			uav_address              : out std_logic_vector(11 downto 0);                    -- address
			uav_burstcount           : out std_logic_vector(2 downto 0);                     -- burstcount
			uav_read                 : out std_logic;                                        -- read
			uav_write                : out std_logic;                                        -- write
			uav_waitrequest          : in  std_logic                     := 'X';             -- waitrequest
			uav_readdatavalid        : in  std_logic                     := 'X';             -- readdatavalid
			uav_byteenable           : out std_logic_vector(3 downto 0);                     -- byteenable
			uav_readdata             : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			uav_writedata            : out std_logic_vector(31 downto 0);                    -- writedata
			uav_lock                 : out std_logic;                                        -- lock
			uav_debugaccess          : out std_logic;                                        -- debugaccess
			av_address               : in  std_logic_vector(9 downto 0)  := (others => 'X'); -- address
			av_waitrequest           : out std_logic;                                        -- waitrequest
			av_byteenable            : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			av_read                  : in  std_logic                     := 'X';             -- read
			av_readdata              : out std_logic_vector(31 downto 0);                    -- readdata
			av_burstcount            : in  std_logic_vector(0 downto 0)  := (others => 'X'); -- burstcount
			av_beginbursttransfer    : in  std_logic                     := 'X';             -- beginbursttransfer
			av_begintransfer         : in  std_logic                     := 'X';             -- begintransfer
			av_chipselect            : in  std_logic                     := 'X';             -- chipselect
			av_readdatavalid         : out std_logic;                                        -- readdatavalid
			av_write                 : in  std_logic                     := 'X';             -- write
			av_writedata             : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			av_lock                  : in  std_logic                     := 'X';             -- lock
			av_debugaccess           : in  std_logic                     := 'X';             -- debugaccess
			uav_clken                : out std_logic;                                        -- clken
			av_clken                 : in  std_logic                     := 'X';             -- clken
			uav_response             : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- response
			av_response              : out std_logic_vector(1 downto 0);                     -- response
			uav_writeresponserequest : out std_logic;                                        -- writeresponserequest
			uav_writeresponsevalid   : in  std_logic                     := 'X';             -- writeresponsevalid
			av_writeresponserequest  : in  std_logic                     := 'X';             -- writeresponserequest
			av_writeresponsevalid    : out std_logic                                         -- writeresponsevalid
		);
	end component fetchmemory_blockram_masterinterface_0_fetchmaster_translator;

	component fetchmemory_blockram_masterinterface_0_memorymaster_translator is
		generic (
			AV_ADDRESS_W                : integer := 32;
			AV_DATA_W                   : integer := 32;
			AV_BURSTCOUNT_W             : integer := 4;
			AV_BYTEENABLE_W             : integer := 4;
			UAV_ADDRESS_W               : integer := 38;
			UAV_BURSTCOUNT_W            : integer := 10;
			USE_READ                    : integer := 1;
			USE_WRITE                   : integer := 1;
			USE_BEGINBURSTTRANSFER      : integer := 0;
			USE_BEGINTRANSFER           : integer := 0;
			USE_CHIPSELECT              : integer := 0;
			USE_BURSTCOUNT              : integer := 1;
			USE_READDATAVALID           : integer := 1;
			USE_WAITREQUEST             : integer := 1;
			USE_READRESPONSE            : integer := 0;
			USE_WRITERESPONSE           : integer := 0;
			AV_SYMBOLS_PER_WORD         : integer := 4;
			AV_ADDRESS_SYMBOLS          : integer := 0;
			AV_BURSTCOUNT_SYMBOLS       : integer := 0;
			AV_CONSTANT_BURST_BEHAVIOR  : integer := 0;
			UAV_CONSTANT_BURST_BEHAVIOR : integer := 0;
			AV_LINEWRAPBURSTS           : integer := 0;
			AV_REGISTERINCOMINGSIGNALS  : integer := 0
		);
		port (
			clk                      : in  std_logic                     := 'X';             -- clk
			reset                    : in  std_logic                     := 'X';             -- reset
			uav_address              : out std_logic_vector(11 downto 0);                    -- address
			uav_burstcount           : out std_logic_vector(2 downto 0);                     -- burstcount
			uav_read                 : out std_logic;                                        -- read
			uav_write                : out std_logic;                                        -- write
			uav_waitrequest          : in  std_logic                     := 'X';             -- waitrequest
			uav_readdatavalid        : in  std_logic                     := 'X';             -- readdatavalid
			uav_byteenable           : out std_logic_vector(3 downto 0);                     -- byteenable
			uav_readdata             : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			uav_writedata            : out std_logic_vector(31 downto 0);                    -- writedata
			uav_lock                 : out std_logic;                                        -- lock
			uav_debugaccess          : out std_logic;                                        -- debugaccess
			av_address               : in  std_logic_vector(9 downto 0)  := (others => 'X'); -- address
			av_waitrequest           : out std_logic;                                        -- waitrequest
			av_byteenable            : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			av_read                  : in  std_logic                     := 'X';             -- read
			av_readdata              : out std_logic_vector(31 downto 0);                    -- readdata
			av_write                 : in  std_logic                     := 'X';             -- write
			av_writedata             : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			av_burstcount            : in  std_logic_vector(0 downto 0)  := (others => 'X'); -- burstcount
			av_beginbursttransfer    : in  std_logic                     := 'X';             -- beginbursttransfer
			av_begintransfer         : in  std_logic                     := 'X';             -- begintransfer
			av_chipselect            : in  std_logic                     := 'X';             -- chipselect
			av_readdatavalid         : out std_logic;                                        -- readdatavalid
			av_lock                  : in  std_logic                     := 'X';             -- lock
			av_debugaccess           : in  std_logic                     := 'X';             -- debugaccess
			uav_clken                : out std_logic;                                        -- clken
			av_clken                 : in  std_logic                     := 'X';             -- clken
			uav_response             : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- response
			av_response              : out std_logic_vector(1 downto 0);                     -- response
			uav_writeresponserequest : out std_logic;                                        -- writeresponserequest
			uav_writeresponsevalid   : in  std_logic                     := 'X';             -- writeresponsevalid
			av_writeresponserequest  : in  std_logic                     := 'X';             -- writeresponserequest
			av_writeresponsevalid    : out std_logic                                         -- writeresponsevalid
		);
	end component fetchmemory_blockram_masterinterface_0_memorymaster_translator;

	signal masterinterface_0_fetchmaster_waitrequest                                         : std_logic;                     -- MasterInterface_0_FetchMaster_translator:av_waitrequest -> MasterInterface_0:fetch_waitrequest
	signal masterinterface_0_fetchmaster_address                                             : std_logic_vector(9 downto 0);  -- MasterInterface_0:fetch_address -> MasterInterface_0_FetchMaster_translator:av_address
	signal masterinterface_0_fetchmaster_read                                                : std_logic;                     -- MasterInterface_0:fetch_read -> MasterInterface_0_FetchMaster_translator:av_read
	signal masterinterface_0_fetchmaster_readdata                                            : std_logic_vector(31 downto 0); -- MasterInterface_0_FetchMaster_translator:av_readdata -> MasterInterface_0:fetch_readdata
	signal masterinterface_0_fetchmaster_byteenable                                          : std_logic_vector(3 downto 0);  -- MasterInterface_0:fetch_byteenable -> MasterInterface_0_FetchMaster_translator:av_byteenable
	signal masterinterface_0_fetchmaster_translator_avalon_universal_master_0_waitrequest    : std_logic;                     -- InstructionMemory_s1_translator:uav_waitrequest -> MasterInterface_0_FetchMaster_translator:uav_waitrequest
	signal masterinterface_0_fetchmaster_translator_avalon_universal_master_0_burstcount     : std_logic_vector(2 downto 0);  -- MasterInterface_0_FetchMaster_translator:uav_burstcount -> InstructionMemory_s1_translator:uav_burstcount
	signal masterinterface_0_fetchmaster_translator_avalon_universal_master_0_writedata      : std_logic_vector(31 downto 0); -- MasterInterface_0_FetchMaster_translator:uav_writedata -> InstructionMemory_s1_translator:uav_writedata
	signal masterinterface_0_fetchmaster_translator_avalon_universal_master_0_address        : std_logic_vector(11 downto 0); -- MasterInterface_0_FetchMaster_translator:uav_address -> InstructionMemory_s1_translator:uav_address
	signal masterinterface_0_fetchmaster_translator_avalon_universal_master_0_lock           : std_logic;                     -- MasterInterface_0_FetchMaster_translator:uav_lock -> InstructionMemory_s1_translator:uav_lock
	signal masterinterface_0_fetchmaster_translator_avalon_universal_master_0_write          : std_logic;                     -- MasterInterface_0_FetchMaster_translator:uav_write -> InstructionMemory_s1_translator:uav_write
	signal masterinterface_0_fetchmaster_translator_avalon_universal_master_0_read           : std_logic;                     -- MasterInterface_0_FetchMaster_translator:uav_read -> InstructionMemory_s1_translator:uav_read
	signal masterinterface_0_fetchmaster_translator_avalon_universal_master_0_readdata       : std_logic_vector(31 downto 0); -- InstructionMemory_s1_translator:uav_readdata -> MasterInterface_0_FetchMaster_translator:uav_readdata
	signal masterinterface_0_fetchmaster_translator_avalon_universal_master_0_debugaccess    : std_logic;                     -- MasterInterface_0_FetchMaster_translator:uav_debugaccess -> InstructionMemory_s1_translator:uav_debugaccess
	signal masterinterface_0_fetchmaster_translator_avalon_universal_master_0_byteenable     : std_logic_vector(3 downto 0);  -- MasterInterface_0_FetchMaster_translator:uav_byteenable -> InstructionMemory_s1_translator:uav_byteenable
	signal masterinterface_0_fetchmaster_translator_avalon_universal_master_0_readdatavalid  : std_logic;                     -- InstructionMemory_s1_translator:uav_readdatavalid -> MasterInterface_0_FetchMaster_translator:uav_readdatavalid
	signal instructionmemory_s1_translator_avalon_anti_slave_0_writedata                     : std_logic_vector(31 downto 0); -- InstructionMemory_s1_translator:av_writedata -> InstructionMemory:writedata
	signal instructionmemory_s1_translator_avalon_anti_slave_0_address                       : std_logic_vector(9 downto 0);  -- InstructionMemory_s1_translator:av_address -> InstructionMemory:address
	signal instructionmemory_s1_translator_avalon_anti_slave_0_chipselect                    : std_logic;                     -- InstructionMemory_s1_translator:av_chipselect -> InstructionMemory:chipselect
	signal instructionmemory_s1_translator_avalon_anti_slave_0_clken                         : std_logic;                     -- InstructionMemory_s1_translator:av_clken -> InstructionMemory:clken
	signal instructionmemory_s1_translator_avalon_anti_slave_0_write                         : std_logic;                     -- InstructionMemory_s1_translator:av_write -> InstructionMemory:write
	signal instructionmemory_s1_translator_avalon_anti_slave_0_readdata                      : std_logic_vector(31 downto 0); -- InstructionMemory:readdata -> InstructionMemory_s1_translator:av_readdata
	signal instructionmemory_s1_translator_avalon_anti_slave_0_debugaccess                   : std_logic;                     -- InstructionMemory_s1_translator:av_debugaccess -> InstructionMemory:debugaccess
	signal instructionmemory_s1_translator_avalon_anti_slave_0_byteenable                    : std_logic_vector(3 downto 0);  -- InstructionMemory_s1_translator:av_byteenable -> InstructionMemory:byteenable
	signal masterinterface_0_memorymaster_waitrequest                                        : std_logic;                     -- MasterInterface_0_MemoryMaster_translator:av_waitrequest -> MasterInterface_0:m_waitrequest
	signal masterinterface_0_memorymaster_writedata                                          : std_logic_vector(31 downto 0); -- MasterInterface_0:m_writedata -> MasterInterface_0_MemoryMaster_translator:av_writedata
	signal masterinterface_0_memorymaster_address                                            : std_logic_vector(9 downto 0);  -- MasterInterface_0:m_address -> MasterInterface_0_MemoryMaster_translator:av_address
	signal masterinterface_0_memorymaster_write                                              : std_logic;                     -- MasterInterface_0:m_write -> MasterInterface_0_MemoryMaster_translator:av_write
	signal masterinterface_0_memorymaster_read                                               : std_logic;                     -- MasterInterface_0:m_read -> MasterInterface_0_MemoryMaster_translator:av_read
	signal masterinterface_0_memorymaster_readdata                                           : std_logic_vector(31 downto 0); -- MasterInterface_0_MemoryMaster_translator:av_readdata -> MasterInterface_0:m_readdata
	signal masterinterface_0_memorymaster_byteenable                                         : std_logic_vector(3 downto 0);  -- MasterInterface_0:m_byteenable -> MasterInterface_0_MemoryMaster_translator:av_byteenable
	signal masterinterface_0_memorymaster_translator_avalon_universal_master_0_waitrequest   : std_logic;                     -- Memory_s1_translator:uav_waitrequest -> MasterInterface_0_MemoryMaster_translator:uav_waitrequest
	signal masterinterface_0_memorymaster_translator_avalon_universal_master_0_burstcount    : std_logic_vector(2 downto 0);  -- MasterInterface_0_MemoryMaster_translator:uav_burstcount -> Memory_s1_translator:uav_burstcount
	signal masterinterface_0_memorymaster_translator_avalon_universal_master_0_writedata     : std_logic_vector(31 downto 0); -- MasterInterface_0_MemoryMaster_translator:uav_writedata -> Memory_s1_translator:uav_writedata
	signal masterinterface_0_memorymaster_translator_avalon_universal_master_0_address       : std_logic_vector(11 downto 0); -- MasterInterface_0_MemoryMaster_translator:uav_address -> Memory_s1_translator:uav_address
	signal masterinterface_0_memorymaster_translator_avalon_universal_master_0_lock          : std_logic;                     -- MasterInterface_0_MemoryMaster_translator:uav_lock -> Memory_s1_translator:uav_lock
	signal masterinterface_0_memorymaster_translator_avalon_universal_master_0_write         : std_logic;                     -- MasterInterface_0_MemoryMaster_translator:uav_write -> Memory_s1_translator:uav_write
	signal masterinterface_0_memorymaster_translator_avalon_universal_master_0_read          : std_logic;                     -- MasterInterface_0_MemoryMaster_translator:uav_read -> Memory_s1_translator:uav_read
	signal masterinterface_0_memorymaster_translator_avalon_universal_master_0_readdata      : std_logic_vector(31 downto 0); -- Memory_s1_translator:uav_readdata -> MasterInterface_0_MemoryMaster_translator:uav_readdata
	signal masterinterface_0_memorymaster_translator_avalon_universal_master_0_debugaccess   : std_logic;                     -- MasterInterface_0_MemoryMaster_translator:uav_debugaccess -> Memory_s1_translator:uav_debugaccess
	signal masterinterface_0_memorymaster_translator_avalon_universal_master_0_byteenable    : std_logic_vector(3 downto 0);  -- MasterInterface_0_MemoryMaster_translator:uav_byteenable -> Memory_s1_translator:uav_byteenable
	signal masterinterface_0_memorymaster_translator_avalon_universal_master_0_readdatavalid : std_logic;                     -- Memory_s1_translator:uav_readdatavalid -> MasterInterface_0_MemoryMaster_translator:uav_readdatavalid
	signal memory_s1_translator_avalon_anti_slave_0_writedata                                : std_logic_vector(31 downto 0); -- Memory_s1_translator:av_writedata -> Memory:writedata
	signal memory_s1_translator_avalon_anti_slave_0_address                                  : std_logic_vector(9 downto 0);  -- Memory_s1_translator:av_address -> Memory:address
	signal memory_s1_translator_avalon_anti_slave_0_chipselect                               : std_logic;                     -- Memory_s1_translator:av_chipselect -> Memory:chipselect
	signal memory_s1_translator_avalon_anti_slave_0_clken                                    : std_logic;                     -- Memory_s1_translator:av_clken -> Memory:clken
	signal memory_s1_translator_avalon_anti_slave_0_write                                    : std_logic;                     -- Memory_s1_translator:av_write -> Memory:write
	signal memory_s1_translator_avalon_anti_slave_0_readdata                                 : std_logic_vector(31 downto 0); -- Memory:readdata -> Memory_s1_translator:av_readdata
	signal memory_s1_translator_avalon_anti_slave_0_byteenable                               : std_logic_vector(3 downto 0);  -- Memory_s1_translator:av_byteenable -> Memory:byteenable
	signal rst_controller_reset_out_reset                                                    : std_logic;                     -- rst_controller:reset_out -> [InstructionMemory:reset, InstructionMemory_s1_translator:reset, MasterInterface_0_FetchMaster_translator:reset, MasterInterface_0_MemoryMaster_translator:reset, Memory:reset, Memory_s1_translator:reset]
	signal rst_controller_reset_out_reset_req                                                : std_logic;                     -- rst_controller:reset_req -> [InstructionMemory:reset_req, Memory:reset_req]
	signal rst_controller_001_reset_out_reset                                                : std_logic;                     -- rst_controller_001:reset_out -> MasterInterface_0:KEY
	signal reset_reset_n_ports_inv                                                           : std_logic;                     -- reset_reset_n:inv -> [rst_controller:reset_in0, rst_controller_001:reset_in0]

begin

	memory : component FetchMemory_Blockram_Memory
		port map (
			clk        => clk_clk,                                             --   clk1.clk
			address    => memory_s1_translator_avalon_anti_slave_0_address,    --     s1.address
			clken      => memory_s1_translator_avalon_anti_slave_0_clken,      --       .clken
			chipselect => memory_s1_translator_avalon_anti_slave_0_chipselect, --       .chipselect
			write      => memory_s1_translator_avalon_anti_slave_0_write,      --       .write
			readdata   => memory_s1_translator_avalon_anti_slave_0_readdata,   --       .readdata
			writedata  => memory_s1_translator_avalon_anti_slave_0_writedata,  --       .writedata
			byteenable => memory_s1_translator_avalon_anti_slave_0_byteenable, --       .byteenable
			reset      => rst_controller_reset_out_reset,                      -- reset1.reset
			reset_req  => rst_controller_reset_out_reset_req                   --       .reset_req
		);

	instructionmemory : component FetchMemory_Blockram_InstructionMemory
		port map (
			clk         => clk_clk,                                                         --   clk1.clk
			address     => instructionmemory_s1_translator_avalon_anti_slave_0_address,     --     s1.address
			debugaccess => instructionmemory_s1_translator_avalon_anti_slave_0_debugaccess, --       .debugaccess
			clken       => instructionmemory_s1_translator_avalon_anti_slave_0_clken,       --       .clken
			chipselect  => instructionmemory_s1_translator_avalon_anti_slave_0_chipselect,  --       .chipselect
			write       => instructionmemory_s1_translator_avalon_anti_slave_0_write,       --       .write
			readdata    => instructionmemory_s1_translator_avalon_anti_slave_0_readdata,    --       .readdata
			writedata   => instructionmemory_s1_translator_avalon_anti_slave_0_writedata,   --       .writedata
			byteenable  => instructionmemory_s1_translator_avalon_anti_slave_0_byteenable,  --       .byteenable
			reset       => rst_controller_reset_out_reset,                                  -- reset1.reset
			reset_req   => rst_controller_reset_out_reset_req                               --       .reset_req
		);

	masterinterface_0 : component RISCV
		port map (
			CLOCK_50          => clk_clk,                                    --   clock_sink.clk
			KEY(0)            => rst_controller_001_reset_out_reset,         --   reset_sink.reset
			fetch_waitrequest => masterinterface_0_fetchmaster_waitrequest,  --  FetchMaster.waitrequest
			fetch_readdata    => masterinterface_0_fetchmaster_readdata,     --             .readdata
			fetch_read        => masterinterface_0_fetchmaster_read,         --             .read
			fetch_address     => masterinterface_0_fetchmaster_address,      --             .address
			fetch_byteenable  => masterinterface_0_fetchmaster_byteenable,   --             .byteenable
			m_waitrequest     => masterinterface_0_memorymaster_waitrequest, -- MemoryMaster.waitrequest
			m_readdata        => masterinterface_0_memorymaster_readdata,    --             .readdata
			m_write           => masterinterface_0_memorymaster_write,       --             .write
			m_read            => masterinterface_0_memorymaster_read,        --             .read
			m_address         => masterinterface_0_memorymaster_address,     --             .address
			m_byteenable      => masterinterface_0_memorymaster_byteenable,  --             .byteenable
			m_writedata       => masterinterface_0_memorymaster_writedata,   --             .writedata
			HEX0              => open,                                       --  conduit_end.export
			HEX1              => open,                                       --             .export
			HEX2              => open,                                       --             .export
			HEX3              => open                                        --             .export
		);

	masterinterface_0_fetchmaster_translator : component fetchmemory_blockram_masterinterface_0_fetchmaster_translator
		generic map (
			AV_ADDRESS_W                => 10,
			AV_DATA_W                   => 32,
			AV_BURSTCOUNT_W             => 1,
			AV_BYTEENABLE_W             => 4,
			UAV_ADDRESS_W               => 12,
			UAV_BURSTCOUNT_W            => 3,
			USE_READ                    => 1,
			USE_WRITE                   => 0,
			USE_BEGINBURSTTRANSFER      => 0,
			USE_BEGINTRANSFER           => 0,
			USE_CHIPSELECT              => 0,
			USE_BURSTCOUNT              => 0,
			USE_READDATAVALID           => 0,
			USE_WAITREQUEST             => 1,
			USE_READRESPONSE            => 0,
			USE_WRITERESPONSE           => 0,
			AV_SYMBOLS_PER_WORD         => 4,
			AV_ADDRESS_SYMBOLS          => 0,
			AV_BURSTCOUNT_SYMBOLS       => 0,
			AV_CONSTANT_BURST_BEHAVIOR  => 0,
			UAV_CONSTANT_BURST_BEHAVIOR => 0,
			AV_LINEWRAPBURSTS           => 0,
			AV_REGISTERINCOMINGSIGNALS  => 0
		)
		port map (
			clk                      => clk_clk,                                                                          --                       clk.clk
			reset                    => rst_controller_reset_out_reset,                                                   --                     reset.reset
			uav_address              => masterinterface_0_fetchmaster_translator_avalon_universal_master_0_address,       -- avalon_universal_master_0.address
			uav_burstcount           => masterinterface_0_fetchmaster_translator_avalon_universal_master_0_burstcount,    --                          .burstcount
			uav_read                 => masterinterface_0_fetchmaster_translator_avalon_universal_master_0_read,          --                          .read
			uav_write                => masterinterface_0_fetchmaster_translator_avalon_universal_master_0_write,         --                          .write
			uav_waitrequest          => masterinterface_0_fetchmaster_translator_avalon_universal_master_0_waitrequest,   --                          .waitrequest
			uav_readdatavalid        => masterinterface_0_fetchmaster_translator_avalon_universal_master_0_readdatavalid, --                          .readdatavalid
			uav_byteenable           => masterinterface_0_fetchmaster_translator_avalon_universal_master_0_byteenable,    --                          .byteenable
			uav_readdata             => masterinterface_0_fetchmaster_translator_avalon_universal_master_0_readdata,      --                          .readdata
			uav_writedata            => masterinterface_0_fetchmaster_translator_avalon_universal_master_0_writedata,     --                          .writedata
			uav_lock                 => masterinterface_0_fetchmaster_translator_avalon_universal_master_0_lock,          --                          .lock
			uav_debugaccess          => masterinterface_0_fetchmaster_translator_avalon_universal_master_0_debugaccess,   --                          .debugaccess
			av_address               => masterinterface_0_fetchmaster_address,                                            --      avalon_anti_master_0.address
			av_waitrequest           => masterinterface_0_fetchmaster_waitrequest,                                        --                          .waitrequest
			av_byteenable            => masterinterface_0_fetchmaster_byteenable,                                         --                          .byteenable
			av_read                  => masterinterface_0_fetchmaster_read,                                               --                          .read
			av_readdata              => masterinterface_0_fetchmaster_readdata,                                           --                          .readdata
			av_burstcount            => "1",                                                                              --               (terminated)
			av_beginbursttransfer    => '0',                                                                              --               (terminated)
			av_begintransfer         => '0',                                                                              --               (terminated)
			av_chipselect            => '0',                                                                              --               (terminated)
			av_readdatavalid         => open,                                                                             --               (terminated)
			av_write                 => '0',                                                                              --               (terminated)
			av_writedata             => "00000000000000000000000000000000",                                               --               (terminated)
			av_lock                  => '0',                                                                              --               (terminated)
			av_debugaccess           => '0',                                                                              --               (terminated)
			uav_clken                => open,                                                                             --               (terminated)
			av_clken                 => '1',                                                                              --               (terminated)
			uav_response             => "00",                                                                             --               (terminated)
			av_response              => open,                                                                             --               (terminated)
			uav_writeresponserequest => open,                                                                             --               (terminated)
			uav_writeresponsevalid   => '0',                                                                              --               (terminated)
			av_writeresponserequest  => '0',                                                                              --               (terminated)
			av_writeresponsevalid    => open                                                                              --               (terminated)
		);

	instructionmemory_s1_translator : component fetchmemory_blockram_instructionmemory_s1_translator
		generic map (
			AV_ADDRESS_W                   => 10,
			AV_DATA_W                      => 32,
			UAV_DATA_W                     => 32,
			AV_BURSTCOUNT_W                => 1,
			AV_BYTEENABLE_W                => 4,
			UAV_BYTEENABLE_W               => 4,
			UAV_ADDRESS_W                  => 12,
			UAV_BURSTCOUNT_W               => 3,
			AV_READLATENCY                 => 1,
			USE_READDATAVALID              => 0,
			USE_WAITREQUEST                => 0,
			USE_UAV_CLKEN                  => 0,
			USE_READRESPONSE               => 0,
			USE_WRITERESPONSE              => 0,
			AV_SYMBOLS_PER_WORD            => 4,
			AV_ADDRESS_SYMBOLS             => 0,
			AV_BURSTCOUNT_SYMBOLS          => 0,
			AV_CONSTANT_BURST_BEHAVIOR     => 0,
			UAV_CONSTANT_BURST_BEHAVIOR    => 0,
			AV_REQUIRE_UNALIGNED_ADDRESSES => 0,
			CHIPSELECT_THROUGH_READLATENCY => 0,
			AV_READ_WAIT_CYCLES            => 0,
			AV_WRITE_WAIT_CYCLES           => 0,
			AV_SETUP_WAIT_CYCLES           => 0,
			AV_DATA_HOLD_CYCLES            => 0
		)
		port map (
			clk                      => clk_clk,                                                                          --                      clk.clk
			reset                    => rst_controller_reset_out_reset,                                                   --                    reset.reset
			uav_address              => masterinterface_0_fetchmaster_translator_avalon_universal_master_0_address,       -- avalon_universal_slave_0.address
			uav_burstcount           => masterinterface_0_fetchmaster_translator_avalon_universal_master_0_burstcount,    --                         .burstcount
			uav_read                 => masterinterface_0_fetchmaster_translator_avalon_universal_master_0_read,          --                         .read
			uav_write                => masterinterface_0_fetchmaster_translator_avalon_universal_master_0_write,         --                         .write
			uav_waitrequest          => masterinterface_0_fetchmaster_translator_avalon_universal_master_0_waitrequest,   --                         .waitrequest
			uav_readdatavalid        => masterinterface_0_fetchmaster_translator_avalon_universal_master_0_readdatavalid, --                         .readdatavalid
			uav_byteenable           => masterinterface_0_fetchmaster_translator_avalon_universal_master_0_byteenable,    --                         .byteenable
			uav_readdata             => masterinterface_0_fetchmaster_translator_avalon_universal_master_0_readdata,      --                         .readdata
			uav_writedata            => masterinterface_0_fetchmaster_translator_avalon_universal_master_0_writedata,     --                         .writedata
			uav_lock                 => masterinterface_0_fetchmaster_translator_avalon_universal_master_0_lock,          --                         .lock
			uav_debugaccess          => masterinterface_0_fetchmaster_translator_avalon_universal_master_0_debugaccess,   --                         .debugaccess
			av_address               => instructionmemory_s1_translator_avalon_anti_slave_0_address,                      --      avalon_anti_slave_0.address
			av_write                 => instructionmemory_s1_translator_avalon_anti_slave_0_write,                        --                         .write
			av_readdata              => instructionmemory_s1_translator_avalon_anti_slave_0_readdata,                     --                         .readdata
			av_writedata             => instructionmemory_s1_translator_avalon_anti_slave_0_writedata,                    --                         .writedata
			av_byteenable            => instructionmemory_s1_translator_avalon_anti_slave_0_byteenable,                   --                         .byteenable
			av_chipselect            => instructionmemory_s1_translator_avalon_anti_slave_0_chipselect,                   --                         .chipselect
			av_clken                 => instructionmemory_s1_translator_avalon_anti_slave_0_clken,                        --                         .clken
			av_debugaccess           => instructionmemory_s1_translator_avalon_anti_slave_0_debugaccess,                  --                         .debugaccess
			av_read                  => open,                                                                             --              (terminated)
			av_begintransfer         => open,                                                                             --              (terminated)
			av_beginbursttransfer    => open,                                                                             --              (terminated)
			av_burstcount            => open,                                                                             --              (terminated)
			av_readdatavalid         => '0',                                                                              --              (terminated)
			av_waitrequest           => '0',                                                                              --              (terminated)
			av_writebyteenable       => open,                                                                             --              (terminated)
			av_lock                  => open,                                                                             --              (terminated)
			uav_clken                => '0',                                                                              --              (terminated)
			av_outputenable          => open,                                                                             --              (terminated)
			uav_response             => open,                                                                             --              (terminated)
			av_response              => "00",                                                                             --              (terminated)
			uav_writeresponserequest => '0',                                                                              --              (terminated)
			uav_writeresponsevalid   => open,                                                                             --              (terminated)
			av_writeresponserequest  => open,                                                                             --              (terminated)
			av_writeresponsevalid    => '0'                                                                               --              (terminated)
		);

	masterinterface_0_memorymaster_translator : component fetchmemory_blockram_masterinterface_0_memorymaster_translator
		generic map (
			AV_ADDRESS_W                => 10,
			AV_DATA_W                   => 32,
			AV_BURSTCOUNT_W             => 1,
			AV_BYTEENABLE_W             => 4,
			UAV_ADDRESS_W               => 12,
			UAV_BURSTCOUNT_W            => 3,
			USE_READ                    => 1,
			USE_WRITE                   => 1,
			USE_BEGINBURSTTRANSFER      => 0,
			USE_BEGINTRANSFER           => 0,
			USE_CHIPSELECT              => 0,
			USE_BURSTCOUNT              => 0,
			USE_READDATAVALID           => 0,
			USE_WAITREQUEST             => 1,
			USE_READRESPONSE            => 0,
			USE_WRITERESPONSE           => 0,
			AV_SYMBOLS_PER_WORD         => 4,
			AV_ADDRESS_SYMBOLS          => 0,
			AV_BURSTCOUNT_SYMBOLS       => 0,
			AV_CONSTANT_BURST_BEHAVIOR  => 0,
			UAV_CONSTANT_BURST_BEHAVIOR => 0,
			AV_LINEWRAPBURSTS           => 0,
			AV_REGISTERINCOMINGSIGNALS  => 0
		)
		port map (
			clk                      => clk_clk,                                                                           --                       clk.clk
			reset                    => rst_controller_reset_out_reset,                                                    --                     reset.reset
			uav_address              => masterinterface_0_memorymaster_translator_avalon_universal_master_0_address,       -- avalon_universal_master_0.address
			uav_burstcount           => masterinterface_0_memorymaster_translator_avalon_universal_master_0_burstcount,    --                          .burstcount
			uav_read                 => masterinterface_0_memorymaster_translator_avalon_universal_master_0_read,          --                          .read
			uav_write                => masterinterface_0_memorymaster_translator_avalon_universal_master_0_write,         --                          .write
			uav_waitrequest          => masterinterface_0_memorymaster_translator_avalon_universal_master_0_waitrequest,   --                          .waitrequest
			uav_readdatavalid        => masterinterface_0_memorymaster_translator_avalon_universal_master_0_readdatavalid, --                          .readdatavalid
			uav_byteenable           => masterinterface_0_memorymaster_translator_avalon_universal_master_0_byteenable,    --                          .byteenable
			uav_readdata             => masterinterface_0_memorymaster_translator_avalon_universal_master_0_readdata,      --                          .readdata
			uav_writedata            => masterinterface_0_memorymaster_translator_avalon_universal_master_0_writedata,     --                          .writedata
			uav_lock                 => masterinterface_0_memorymaster_translator_avalon_universal_master_0_lock,          --                          .lock
			uav_debugaccess          => masterinterface_0_memorymaster_translator_avalon_universal_master_0_debugaccess,   --                          .debugaccess
			av_address               => masterinterface_0_memorymaster_address,                                            --      avalon_anti_master_0.address
			av_waitrequest           => masterinterface_0_memorymaster_waitrequest,                                        --                          .waitrequest
			av_byteenable            => masterinterface_0_memorymaster_byteenable,                                         --                          .byteenable
			av_read                  => masterinterface_0_memorymaster_read,                                               --                          .read
			av_readdata              => masterinterface_0_memorymaster_readdata,                                           --                          .readdata
			av_write                 => masterinterface_0_memorymaster_write,                                              --                          .write
			av_writedata             => masterinterface_0_memorymaster_writedata,                                          --                          .writedata
			av_burstcount            => "1",                                                                               --               (terminated)
			av_beginbursttransfer    => '0',                                                                               --               (terminated)
			av_begintransfer         => '0',                                                                               --               (terminated)
			av_chipselect            => '0',                                                                               --               (terminated)
			av_readdatavalid         => open,                                                                              --               (terminated)
			av_lock                  => '0',                                                                               --               (terminated)
			av_debugaccess           => '0',                                                                               --               (terminated)
			uav_clken                => open,                                                                              --               (terminated)
			av_clken                 => '1',                                                                               --               (terminated)
			uav_response             => "00",                                                                              --               (terminated)
			av_response              => open,                                                                              --               (terminated)
			uav_writeresponserequest => open,                                                                              --               (terminated)
			uav_writeresponsevalid   => '0',                                                                               --               (terminated)
			av_writeresponserequest  => '0',                                                                               --               (terminated)
			av_writeresponsevalid    => open                                                                               --               (terminated)
		);

	memory_s1_translator : component fetchmemory_blockram_memory_s1_translator
		generic map (
			AV_ADDRESS_W                   => 10,
			AV_DATA_W                      => 32,
			UAV_DATA_W                     => 32,
			AV_BURSTCOUNT_W                => 1,
			AV_BYTEENABLE_W                => 4,
			UAV_BYTEENABLE_W               => 4,
			UAV_ADDRESS_W                  => 12,
			UAV_BURSTCOUNT_W               => 3,
			AV_READLATENCY                 => 1,
			USE_READDATAVALID              => 0,
			USE_WAITREQUEST                => 0,
			USE_UAV_CLKEN                  => 0,
			USE_READRESPONSE               => 0,
			USE_WRITERESPONSE              => 0,
			AV_SYMBOLS_PER_WORD            => 4,
			AV_ADDRESS_SYMBOLS             => 0,
			AV_BURSTCOUNT_SYMBOLS          => 0,
			AV_CONSTANT_BURST_BEHAVIOR     => 0,
			UAV_CONSTANT_BURST_BEHAVIOR    => 0,
			AV_REQUIRE_UNALIGNED_ADDRESSES => 0,
			CHIPSELECT_THROUGH_READLATENCY => 0,
			AV_READ_WAIT_CYCLES            => 0,
			AV_WRITE_WAIT_CYCLES           => 0,
			AV_SETUP_WAIT_CYCLES           => 0,
			AV_DATA_HOLD_CYCLES            => 0
		)
		port map (
			clk                      => clk_clk,                                                                           --                      clk.clk
			reset                    => rst_controller_reset_out_reset,                                                    --                    reset.reset
			uav_address              => masterinterface_0_memorymaster_translator_avalon_universal_master_0_address,       -- avalon_universal_slave_0.address
			uav_burstcount           => masterinterface_0_memorymaster_translator_avalon_universal_master_0_burstcount,    --                         .burstcount
			uav_read                 => masterinterface_0_memorymaster_translator_avalon_universal_master_0_read,          --                         .read
			uav_write                => masterinterface_0_memorymaster_translator_avalon_universal_master_0_write,         --                         .write
			uav_waitrequest          => masterinterface_0_memorymaster_translator_avalon_universal_master_0_waitrequest,   --                         .waitrequest
			uav_readdatavalid        => masterinterface_0_memorymaster_translator_avalon_universal_master_0_readdatavalid, --                         .readdatavalid
			uav_byteenable           => masterinterface_0_memorymaster_translator_avalon_universal_master_0_byteenable,    --                         .byteenable
			uav_readdata             => masterinterface_0_memorymaster_translator_avalon_universal_master_0_readdata,      --                         .readdata
			uav_writedata            => masterinterface_0_memorymaster_translator_avalon_universal_master_0_writedata,     --                         .writedata
			uav_lock                 => masterinterface_0_memorymaster_translator_avalon_universal_master_0_lock,          --                         .lock
			uav_debugaccess          => masterinterface_0_memorymaster_translator_avalon_universal_master_0_debugaccess,   --                         .debugaccess
			av_address               => memory_s1_translator_avalon_anti_slave_0_address,                                  --      avalon_anti_slave_0.address
			av_write                 => memory_s1_translator_avalon_anti_slave_0_write,                                    --                         .write
			av_readdata              => memory_s1_translator_avalon_anti_slave_0_readdata,                                 --                         .readdata
			av_writedata             => memory_s1_translator_avalon_anti_slave_0_writedata,                                --                         .writedata
			av_byteenable            => memory_s1_translator_avalon_anti_slave_0_byteenable,                               --                         .byteenable
			av_chipselect            => memory_s1_translator_avalon_anti_slave_0_chipselect,                               --                         .chipselect
			av_clken                 => memory_s1_translator_avalon_anti_slave_0_clken,                                    --                         .clken
			av_read                  => open,                                                                              --              (terminated)
			av_begintransfer         => open,                                                                              --              (terminated)
			av_beginbursttransfer    => open,                                                                              --              (terminated)
			av_burstcount            => open,                                                                              --              (terminated)
			av_readdatavalid         => '0',                                                                               --              (terminated)
			av_waitrequest           => '0',                                                                               --              (terminated)
			av_writebyteenable       => open,                                                                              --              (terminated)
			av_lock                  => open,                                                                              --              (terminated)
			uav_clken                => '0',                                                                               --              (terminated)
			av_debugaccess           => open,                                                                              --              (terminated)
			av_outputenable          => open,                                                                              --              (terminated)
			uav_response             => open,                                                                              --              (terminated)
			av_response              => "00",                                                                              --              (terminated)
			uav_writeresponserequest => '0',                                                                               --              (terminated)
			uav_writeresponsevalid   => open,                                                                              --              (terminated)
			av_writeresponserequest  => open,                                                                              --              (terminated)
			av_writeresponsevalid    => '0'                                                                                --              (terminated)
		);

	rst_controller : component fetchmemory_blockram_rst_controller
		generic map (
			NUM_RESET_INPUTS        => 1,
			OUTPUT_RESET_SYNC_EDGES => "deassert",
			SYNC_DEPTH              => 2,
			RESET_REQUEST_PRESENT   => 1
		)
		port map (
			reset_in0  => reset_reset_n_ports_inv,            -- reset_in0.reset
			clk        => clk_clk,                            --       clk.clk
			reset_out  => rst_controller_reset_out_reset,     -- reset_out.reset
			reset_req  => rst_controller_reset_out_reset_req, --          .reset_req
			reset_in1  => '0',                                -- (terminated)
			reset_in2  => '0',                                -- (terminated)
			reset_in3  => '0',                                -- (terminated)
			reset_in4  => '0',                                -- (terminated)
			reset_in5  => '0',                                -- (terminated)
			reset_in6  => '0',                                -- (terminated)
			reset_in7  => '0',                                -- (terminated)
			reset_in8  => '0',                                -- (terminated)
			reset_in9  => '0',                                -- (terminated)
			reset_in10 => '0',                                -- (terminated)
			reset_in11 => '0',                                -- (terminated)
			reset_in12 => '0',                                -- (terminated)
			reset_in13 => '0',                                -- (terminated)
			reset_in14 => '0',                                -- (terminated)
			reset_in15 => '0'                                 -- (terminated)
		);

	rst_controller_001 : component fetchmemory_blockram_rst_controller_001
		generic map (
			NUM_RESET_INPUTS        => 1,
			OUTPUT_RESET_SYNC_EDGES => "both",
			SYNC_DEPTH              => 2,
			RESET_REQUEST_PRESENT   => 0
		)
		port map (
			reset_in0  => reset_reset_n_ports_inv,            -- reset_in0.reset
			clk        => clk_clk,                            --       clk.clk
			reset_out  => rst_controller_001_reset_out_reset, -- reset_out.reset
			reset_req  => open,                               -- (terminated)
			reset_in1  => '0',                                -- (terminated)
			reset_in2  => '0',                                -- (terminated)
			reset_in3  => '0',                                -- (terminated)
			reset_in4  => '0',                                -- (terminated)
			reset_in5  => '0',                                -- (terminated)
			reset_in6  => '0',                                -- (terminated)
			reset_in7  => '0',                                -- (terminated)
			reset_in8  => '0',                                -- (terminated)
			reset_in9  => '0',                                -- (terminated)
			reset_in10 => '0',                                -- (terminated)
			reset_in11 => '0',                                -- (terminated)
			reset_in12 => '0',                                -- (terminated)
			reset_in13 => '0',                                -- (terminated)
			reset_in14 => '0',                                -- (terminated)
			reset_in15 => '0'                                 -- (terminated)
		);

	reset_reset_n_ports_inv <= not reset_reset_n;

end architecture rtl; -- of FetchMemory_Blockram
