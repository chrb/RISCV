-- SDRAM_tb.vhd

-- Generated using ACDS version 13.0sp1 232 at 2016.02.05.11:39:02

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity SDRAM_tb is
end entity SDRAM_tb;

architecture rtl of SDRAM_tb is
	component SDRAM is
		port (
			clk_clk       : in std_logic := 'X'; -- clk
			reset_reset_n : in std_logic := 'X'  -- reset_n
		);
	end component SDRAM;

	component altera_avalon_clock_source is
		generic (
			CLOCK_RATE : positive := 10;
			CLOCK_UNIT : positive := 1000000
		);
		port (
			clk : out std_logic   -- clk
		);
	end component altera_avalon_clock_source;

	component altera_avalon_reset_source is
		generic (
			ASSERT_HIGH_RESET    : integer := 1;
			INITIAL_RESET_CYCLES : integer := 0
		);
		port (
			reset : out std_logic;        -- reset_n
			clk   : in  std_logic := 'X'  -- clk
		);
	end component altera_avalon_reset_source;

	signal sdram_inst_clk_bfm_clk_clk       : std_logic; -- SDRAM_inst_clk_bfm:clk -> [SDRAM_inst:clk_clk, SDRAM_inst_reset_bfm:clk]
	signal sdram_inst_reset_bfm_reset_reset : std_logic; -- SDRAM_inst_reset_bfm:reset -> SDRAM_inst:reset_reset_n

begin

	sdram_inst : component SDRAM
		port map (
			clk_clk       => sdram_inst_clk_bfm_clk_clk,       --   clk.clk
			reset_reset_n => sdram_inst_reset_bfm_reset_reset  -- reset.reset_n
		);

	sdram_inst_clk_bfm : component altera_avalon_clock_source
		generic map (
			CLOCK_RATE => 50000000,
			CLOCK_UNIT => 1
		)
		port map (
			clk => sdram_inst_clk_bfm_clk_clk  -- clk.clk
		);

	sdram_inst_reset_bfm : component altera_avalon_reset_source
		generic map (
			ASSERT_HIGH_RESET    => 0,
			INITIAL_RESET_CYCLES => 50
		)
		port map (
			reset => sdram_inst_reset_bfm_reset_reset, -- reset.reset_n
			clk   => sdram_inst_clk_bfm_clk_clk        --   clk.clk
		);

end architecture rtl; -- of SDRAM_tb
